module dataMemory(clock, memWrite, address, dataIn, out);
	input clock, memWrite;
	input [31:0] dataIn;
	input[14:0] address;
	output [127:0] out;
	wire [14:0]x;

	reg[31:0] word[32 * 1024 - 1:0];  //32767

	
	always @(posedge clock) begin
		if (memWrite)begin
			word[address] <= dataIn;
		end
	end
	assign out = {word[address + 15'd3], word[address + 15'd2], word[address + 15'd1], word[address]};
	assign x = address + 15'd3;

	always @(clock)begin
		
		word[15'd1024] <= 32'd100;
		word[15'd1025] <= 32'd101;
		word[15'd1026] <= 32'd102;
		word[15'd1027] <= 32'd103;
		word[15'd1028] <= 32'd104;
		word[15'd1029] <= 32'd105;
		word[15'd1030] <= 32'd106;
		word[15'd1031] <= 32'd107;
		word[15'd1032] <= 32'd108;
		word[15'd1033] <= 32'd109;
		word[15'd1034] <= 32'd110;
		word[15'd1035] <= 32'd111;
		word[15'd1036] <= 32'd112;
		word[15'd1037] <= 32'd113;
		word[15'd1038] <= 32'd114;
		word[15'd1039] <= 32'd115;
		word[15'd1040] <= 32'd116;
		word[15'd1041] <= 32'd117;
		word[15'd1042] <= 32'd118;
		word[15'd1043] <= 32'd119;
		word[15'd1044] <= 32'd120;
		word[15'd1045] <= 32'd121;
		word[15'd1046] <= 32'd122;
		word[15'd1047] <= 32'd123;
		word[15'd1048] <= 32'd124;
		word[15'd1049] <= 32'd125;
		word[15'd1050] <= 32'd126;
		word[15'd1051] <= 32'd127;
		word[15'd1052] <= 32'd128;
		word[15'd1053] <= 32'd129;
		word[15'd1054] <= 32'd130;
		word[15'd1055] <= 32'd131;
		word[15'd1056] <= 32'd132;
		word[15'd1057] <= 32'd133;
		word[15'd1058] <= 32'd134;
		word[15'd1059] <= 32'd135;
		word[15'd1060] <= 32'd136;
		word[15'd1061] <= 32'd137;
		word[15'd1062] <= 32'd138;
		word[15'd1063] <= 32'd139;
		word[15'd1064] <= 32'd140;
		word[15'd1065] <= 32'd141;
		word[15'd1066] <= 32'd142;
		word[15'd1067] <= 32'd143;
		word[15'd1068] <= 32'd144;
		word[15'd1069] <= 32'd145;
		word[15'd1070] <= 32'd146;
		word[15'd1071] <= 32'd147;
		word[15'd1072] <= 32'd148;
		word[15'd1073] <= 32'd149;
		word[15'd1074] <= 32'd150;
		word[15'd1075] <= 32'd151;
		word[15'd1076] <= 32'd152;
		word[15'd1077] <= 32'd153;
		word[15'd1078] <= 32'd154;
		word[15'd1079] <= 32'd155;
		word[15'd1080] <= 32'd156;
		word[15'd1081] <= 32'd157;
		word[15'd1082] <= 32'd158;
		word[15'd1083] <= 32'd159;
		word[15'd1084] <= 32'd160;
		word[15'd1085] <= 32'd161;
		word[15'd1086] <= 32'd162;
		word[15'd1087] <= 32'd163;
		word[15'd1088] <= 32'd164;
		word[15'd1089] <= 32'd165;
		word[15'd1090] <= 32'd166;
		word[15'd1091] <= 32'd167;
		word[15'd1092] <= 32'd168;
		word[15'd1093] <= 32'd169;
		word[15'd1094] <= 32'd170;
		word[15'd1095] <= 32'd171;
		word[15'd1096] <= 32'd172;
		word[15'd1097] <= 32'd173;
		word[15'd1098] <= 32'd174;
		word[15'd1099] <= 32'd175;
		word[15'd1100] <= 32'd176;
		word[15'd1101] <= 32'd177;
		word[15'd1102] <= 32'd178;
		word[15'd1103] <= 32'd179;
		word[15'd1104] <= 32'd180;
		word[15'd1105] <= 32'd181;
		word[15'd1106] <= 32'd182;
		word[15'd1107] <= 32'd183;
		word[15'd1108] <= 32'd184;
		word[15'd1109] <= 32'd185;
		word[15'd1110] <= 32'd186;
		word[15'd1111] <= 32'd187;
		word[15'd1112] <= 32'd188;
		word[15'd1113] <= 32'd189;
		word[15'd1114] <= 32'd190;
		word[15'd1115] <= 32'd191;
		word[15'd1116] <= 32'd192;
		word[15'd1117] <= 32'd193;
		word[15'd1118] <= 32'd194;
		word[15'd1119] <= 32'd195;
		word[15'd1120] <= 32'd196;
		word[15'd1121] <= 32'd197;
		word[15'd1122] <= 32'd198;
		word[15'd1123] <= 32'd199;
		word[15'd1124] <= 32'd200;
		word[15'd1125] <= 32'd201;
		word[15'd1126] <= 32'd202;
		word[15'd1127] <= 32'd203;
		word[15'd1128] <= 32'd204;
		word[15'd1129] <= 32'd205;
		word[15'd1130] <= 32'd206;
		word[15'd1131] <= 32'd207;
		word[15'd1132] <= 32'd208;
		word[15'd1133] <= 32'd209;
		word[15'd1134] <= 32'd210;
		word[15'd1135] <= 32'd211;
		word[15'd1136] <= 32'd212;
		word[15'd1137] <= 32'd213;
		word[15'd1138] <= 32'd214;
		word[15'd1139] <= 32'd215;
		word[15'd1140] <= 32'd216;
		word[15'd1141] <= 32'd217;
		word[15'd1142] <= 32'd218;
		word[15'd1143] <= 32'd219;
		word[15'd1144] <= 32'd220;
		word[15'd1145] <= 32'd221;
		word[15'd1146] <= 32'd222;
		word[15'd1147] <= 32'd223;
		word[15'd1148] <= 32'd224;
		word[15'd1149] <= 32'd225;
		word[15'd1150] <= 32'd226;
		word[15'd1151] <= 32'd227;
		word[15'd1152] <= 32'd228;
		word[15'd1153] <= 32'd229;
		word[15'd1154] <= 32'd230;
		word[15'd1155] <= 32'd231;
		word[15'd1156] <= 32'd232;
		word[15'd1157] <= 32'd233;
		word[15'd1158] <= 32'd234;
		word[15'd1159] <= 32'd235;
		word[15'd1160] <= 32'd236;
		word[15'd1161] <= 32'd237;
		word[15'd1162] <= 32'd238;
		word[15'd1163] <= 32'd239;
		word[15'd1164] <= 32'd240;
		word[15'd1165] <= 32'd241;
		word[15'd1166] <= 32'd242;
		word[15'd1167] <= 32'd243;
		word[15'd1168] <= 32'd244;
		word[15'd1169] <= 32'd245;
		word[15'd1170] <= 32'd246;
		word[15'd1171] <= 32'd247;
		word[15'd1172] <= 32'd248;
		word[15'd1173] <= 32'd249;
		word[15'd1174] <= 32'd250;
		word[15'd1175] <= 32'd251;
		word[15'd1176] <= 32'd252;
		word[15'd1177] <= 32'd253;
		word[15'd1178] <= 32'd254;
		word[15'd1179] <= 32'd255;
		word[15'd1180] <= 32'd256;
		word[15'd1181] <= 32'd257;
		word[15'd1182] <= 32'd258;
		word[15'd1183] <= 32'd259;
		word[15'd1184] <= 32'd260;
		word[15'd1185] <= 32'd261;
		word[15'd1186] <= 32'd262;
		word[15'd1187] <= 32'd263;
		word[15'd1188] <= 32'd264;
		word[15'd1189] <= 32'd265;
		word[15'd1190] <= 32'd266;
		word[15'd1191] <= 32'd267;
		word[15'd1192] <= 32'd268;
		word[15'd1193] <= 32'd269;
		word[15'd1194] <= 32'd270;
		word[15'd1195] <= 32'd271;
		word[15'd1196] <= 32'd272;
		word[15'd1197] <= 32'd273;
		word[15'd1198] <= 32'd274;
		word[15'd1199] <= 32'd275;
		word[15'd1200] <= 32'd276;
		word[15'd1201] <= 32'd277;
		word[15'd1202] <= 32'd278;
		word[15'd1203] <= 32'd279;
		word[15'd1204] <= 32'd280;
		word[15'd1205] <= 32'd281;
		word[15'd1206] <= 32'd282;
		word[15'd1207] <= 32'd283;
		word[15'd1208] <= 32'd284;
		word[15'd1209] <= 32'd285;
		word[15'd1210] <= 32'd286;
		word[15'd1211] <= 32'd287;
		word[15'd1212] <= 32'd288;
		word[15'd1213] <= 32'd289;
		word[15'd1214] <= 32'd290;
		word[15'd1215] <= 32'd291;
		word[15'd1216] <= 32'd292;
		word[15'd1217] <= 32'd293;
		word[15'd1218] <= 32'd294;
		word[15'd1219] <= 32'd295;
		word[15'd1220] <= 32'd296;
		word[15'd1221] <= 32'd297;
		word[15'd1222] <= 32'd298;
		word[15'd1223] <= 32'd299;
		word[15'd1224] <= 32'd300;
		word[15'd1225] <= 32'd301;
		word[15'd1226] <= 32'd302;
		word[15'd1227] <= 32'd303;
		word[15'd1228] <= 32'd304;
		word[15'd1229] <= 32'd305;
		word[15'd1230] <= 32'd306;
		word[15'd1231] <= 32'd307;
		word[15'd1232] <= 32'd308;
		word[15'd1233] <= 32'd309;
		word[15'd1234] <= 32'd310;
		word[15'd1235] <= 32'd311;
		word[15'd1236] <= 32'd312;
		word[15'd1237] <= 32'd313;
		word[15'd1238] <= 32'd314;
		word[15'd1239] <= 32'd315;
		word[15'd1240] <= 32'd316;
		word[15'd1241] <= 32'd317;
		word[15'd1242] <= 32'd318;
		word[15'd1243] <= 32'd319;
		word[15'd1244] <= 32'd320;
		word[15'd1245] <= 32'd321;
		word[15'd1246] <= 32'd322;
		word[15'd1247] <= 32'd323;
		word[15'd1248] <= 32'd324;
		word[15'd1249] <= 32'd325;
		word[15'd1250] <= 32'd326;
		word[15'd1251] <= 32'd327;
		word[15'd1252] <= 32'd328;
		word[15'd1253] <= 32'd329;
		word[15'd1254] <= 32'd330;
		word[15'd1255] <= 32'd331;
		word[15'd1256] <= 32'd332;
		word[15'd1257] <= 32'd333;
		word[15'd1258] <= 32'd334;
		word[15'd1259] <= 32'd335;
		word[15'd1260] <= 32'd336;
		word[15'd1261] <= 32'd337;
		word[15'd1262] <= 32'd338;
		word[15'd1263] <= 32'd339;
		word[15'd1264] <= 32'd340;
		word[15'd1265] <= 32'd341;
		word[15'd1266] <= 32'd342;
		word[15'd1267] <= 32'd343;
		word[15'd1268] <= 32'd344;
		word[15'd1269] <= 32'd345;
		word[15'd1270] <= 32'd346;
		word[15'd1271] <= 32'd347;
		word[15'd1272] <= 32'd348;
		word[15'd1273] <= 32'd349;
		word[15'd1274] <= 32'd350;
		word[15'd1275] <= 32'd351;
		word[15'd1276] <= 32'd352;
		word[15'd1277] <= 32'd353;
		word[15'd1278] <= 32'd354;
		word[15'd1279] <= 32'd355;
		word[15'd1280] <= 32'd356;
		word[15'd1281] <= 32'd357;
		word[15'd1282] <= 32'd358;
		word[15'd1283] <= 32'd359;
		word[15'd1284] <= 32'd360;
		word[15'd1285] <= 32'd361;
		word[15'd1286] <= 32'd362;
		word[15'd1287] <= 32'd363;
		word[15'd1288] <= 32'd364;
		word[15'd1289] <= 32'd365;
		word[15'd1290] <= 32'd366;
		word[15'd1291] <= 32'd367;
		word[15'd1292] <= 32'd368;
		word[15'd1293] <= 32'd369;
		word[15'd1294] <= 32'd370;
		word[15'd1295] <= 32'd371;
		word[15'd1296] <= 32'd372;
		word[15'd1297] <= 32'd373;
		word[15'd1298] <= 32'd374;
		word[15'd1299] <= 32'd375;
		word[15'd1300] <= 32'd376;
		word[15'd1301] <= 32'd377;
		word[15'd1302] <= 32'd378;
		word[15'd1303] <= 32'd379;
		word[15'd1304] <= 32'd380;
		word[15'd1305] <= 32'd381;
		word[15'd1306] <= 32'd382;
		word[15'd1307] <= 32'd383;
		word[15'd1308] <= 32'd384;
		word[15'd1309] <= 32'd385;
		word[15'd1310] <= 32'd386;
		word[15'd1311] <= 32'd387;
		word[15'd1312] <= 32'd388;
		word[15'd1313] <= 32'd389;
		word[15'd1314] <= 32'd390;
		word[15'd1315] <= 32'd391;
		word[15'd1316] <= 32'd392;
		word[15'd1317] <= 32'd393;
		word[15'd1318] <= 32'd394;
		word[15'd1319] <= 32'd395;
		word[15'd1320] <= 32'd396;
		word[15'd1321] <= 32'd397;
		word[15'd1322] <= 32'd398;
		word[15'd1323] <= 32'd399;
		word[15'd1324] <= 32'd400;
		word[15'd1325] <= 32'd401;
		word[15'd1326] <= 32'd402;
		word[15'd1327] <= 32'd403;
		word[15'd1328] <= 32'd404;
		word[15'd1329] <= 32'd405;
		word[15'd1330] <= 32'd406;
		word[15'd1331] <= 32'd407;
		word[15'd1332] <= 32'd408;
		word[15'd1333] <= 32'd409;
		word[15'd1334] <= 32'd410;
		word[15'd1335] <= 32'd411;
		word[15'd1336] <= 32'd412;
		word[15'd1337] <= 32'd413;
		word[15'd1338] <= 32'd414;
		word[15'd1339] <= 32'd415;
		word[15'd1340] <= 32'd416;
		word[15'd1341] <= 32'd417;
		word[15'd1342] <= 32'd418;
		word[15'd1343] <= 32'd419;
		word[15'd1344] <= 32'd420;
		word[15'd1345] <= 32'd421;
		word[15'd1346] <= 32'd422;
		word[15'd1347] <= 32'd423;
		word[15'd1348] <= 32'd424;
		word[15'd1349] <= 32'd425;
		word[15'd1350] <= 32'd426;
		word[15'd1351] <= 32'd427;
		word[15'd1352] <= 32'd428;
		word[15'd1353] <= 32'd429;
		word[15'd1354] <= 32'd430;
		word[15'd1355] <= 32'd431;
		word[15'd1356] <= 32'd432;
		word[15'd1357] <= 32'd433;
		word[15'd1358] <= 32'd434;
		word[15'd1359] <= 32'd435;
		word[15'd1360] <= 32'd436;
		word[15'd1361] <= 32'd437;
		word[15'd1362] <= 32'd438;
		word[15'd1363] <= 32'd439;
		word[15'd1364] <= 32'd440;
		word[15'd1365] <= 32'd441;
		word[15'd1366] <= 32'd442;
		word[15'd1367] <= 32'd443;
		word[15'd1368] <= 32'd444;
		word[15'd1369] <= 32'd445;
		word[15'd1370] <= 32'd446;
		word[15'd1371] <= 32'd447;
		word[15'd1372] <= 32'd448;
		word[15'd1373] <= 32'd449;
		word[15'd1374] <= 32'd450;
		word[15'd1375] <= 32'd451;
		word[15'd1376] <= 32'd452;
		word[15'd1377] <= 32'd453;
		word[15'd1378] <= 32'd454;
		word[15'd1379] <= 32'd455;
		word[15'd1380] <= 32'd456;
		word[15'd1381] <= 32'd457;
		word[15'd1382] <= 32'd458;
		word[15'd1383] <= 32'd459;
		word[15'd1384] <= 32'd460;
		word[15'd1385] <= 32'd461;
		word[15'd1386] <= 32'd462;
		word[15'd1387] <= 32'd463;
		word[15'd1388] <= 32'd464;
		word[15'd1389] <= 32'd465;
		word[15'd1390] <= 32'd466;
		word[15'd1391] <= 32'd467;
		word[15'd1392] <= 32'd468;
		word[15'd1393] <= 32'd469;
		word[15'd1394] <= 32'd470;
		word[15'd1395] <= 32'd471;
		word[15'd1396] <= 32'd472;
		word[15'd1397] <= 32'd473;
		word[15'd1398] <= 32'd474;
		word[15'd1399] <= 32'd475;
		word[15'd1400] <= 32'd476;
		word[15'd1401] <= 32'd477;
		word[15'd1402] <= 32'd478;
		word[15'd1403] <= 32'd479;
		word[15'd1404] <= 32'd480;
		word[15'd1405] <= 32'd481;
		word[15'd1406] <= 32'd482;
		word[15'd1407] <= 32'd483;
		word[15'd1408] <= 32'd484;
		word[15'd1409] <= 32'd485;
		word[15'd1410] <= 32'd486;
		word[15'd1411] <= 32'd487;
		word[15'd1412] <= 32'd488;
		word[15'd1413] <= 32'd489;
		word[15'd1414] <= 32'd490;
		word[15'd1415] <= 32'd491;
		word[15'd1416] <= 32'd492;
		word[15'd1417] <= 32'd493;
		word[15'd1418] <= 32'd494;
		word[15'd1419] <= 32'd495;
		word[15'd1420] <= 32'd496;
		word[15'd1421] <= 32'd497;
		word[15'd1422] <= 32'd498;
		word[15'd1423] <= 32'd499;
		word[15'd1424] <= 32'd500;
		word[15'd1425] <= 32'd501;
		word[15'd1426] <= 32'd502;
		word[15'd1427] <= 32'd503;
		word[15'd1428] <= 32'd504;
		word[15'd1429] <= 32'd505;
		word[15'd1430] <= 32'd506;
		word[15'd1431] <= 32'd507;
		word[15'd1432] <= 32'd508;
		word[15'd1433] <= 32'd509;
		word[15'd1434] <= 32'd510;
		word[15'd1435] <= 32'd511;
		word[15'd1436] <= 32'd512;
		word[15'd1437] <= 32'd513;
		word[15'd1438] <= 32'd514;
		word[15'd1439] <= 32'd515;
		word[15'd1440] <= 32'd516;
		word[15'd1441] <= 32'd517;
		word[15'd1442] <= 32'd518;
		word[15'd1443] <= 32'd519;
		word[15'd1444] <= 32'd520;
		word[15'd1445] <= 32'd521;
		word[15'd1446] <= 32'd522;
		word[15'd1447] <= 32'd523;
		word[15'd1448] <= 32'd524;
		word[15'd1449] <= 32'd525;
		word[15'd1450] <= 32'd526;
		word[15'd1451] <= 32'd527;
		word[15'd1452] <= 32'd528;
		word[15'd1453] <= 32'd529;
		word[15'd1454] <= 32'd530;
		word[15'd1455] <= 32'd531;
		word[15'd1456] <= 32'd532;
		word[15'd1457] <= 32'd533;
		word[15'd1458] <= 32'd534;
		word[15'd1459] <= 32'd535;
		word[15'd1460] <= 32'd536;
		word[15'd1461] <= 32'd537;
		word[15'd1462] <= 32'd538;
		word[15'd1463] <= 32'd539;
		word[15'd1464] <= 32'd540;
		word[15'd1465] <= 32'd541;
		word[15'd1466] <= 32'd542;
		word[15'd1467] <= 32'd543;
		word[15'd1468] <= 32'd544;
		word[15'd1469] <= 32'd545;
		word[15'd1470] <= 32'd546;
		word[15'd1471] <= 32'd547;
		word[15'd1472] <= 32'd548;
		word[15'd1473] <= 32'd549;
		word[15'd1474] <= 32'd550;
		word[15'd1475] <= 32'd551;
		word[15'd1476] <= 32'd552;
		word[15'd1477] <= 32'd553;
		word[15'd1478] <= 32'd554;
		word[15'd1479] <= 32'd555;
		word[15'd1480] <= 32'd556;
		word[15'd1481] <= 32'd557;
		word[15'd1482] <= 32'd558;
		word[15'd1483] <= 32'd559;
		word[15'd1484] <= 32'd560;
		word[15'd1485] <= 32'd561;
		word[15'd1486] <= 32'd562;
		word[15'd1487] <= 32'd563;
		word[15'd1488] <= 32'd564;
		word[15'd1489] <= 32'd565;
		word[15'd1490] <= 32'd566;
		word[15'd1491] <= 32'd567;
		word[15'd1492] <= 32'd568;
		word[15'd1493] <= 32'd569;
		word[15'd1494] <= 32'd570;
		word[15'd1495] <= 32'd571;
		word[15'd1496] <= 32'd572;
		word[15'd1497] <= 32'd573;
		word[15'd1498] <= 32'd574;
		word[15'd1499] <= 32'd575;
		word[15'd1500] <= 32'd576;
		word[15'd1501] <= 32'd577;
		word[15'd1502] <= 32'd578;
		word[15'd1503] <= 32'd579;
		word[15'd1504] <= 32'd580;
		word[15'd1505] <= 32'd581;
		word[15'd1506] <= 32'd582;
		word[15'd1507] <= 32'd583;
		word[15'd1508] <= 32'd584;
		word[15'd1509] <= 32'd585;
		word[15'd1510] <= 32'd586;
		word[15'd1511] <= 32'd587;
		word[15'd1512] <= 32'd588;
		word[15'd1513] <= 32'd589;
		word[15'd1514] <= 32'd590;
		word[15'd1515] <= 32'd591;
		word[15'd1516] <= 32'd592;
		word[15'd1517] <= 32'd593;
		word[15'd1518] <= 32'd594;
		word[15'd1519] <= 32'd595;
		word[15'd1520] <= 32'd596;
		word[15'd1521] <= 32'd597;
		word[15'd1522] <= 32'd598;
		word[15'd1523] <= 32'd599;
		word[15'd1524] <= 32'd600;
		word[15'd1525] <= 32'd601;
		word[15'd1526] <= 32'd602;
		word[15'd1527] <= 32'd603;
		word[15'd1528] <= 32'd604;
		word[15'd1529] <= 32'd605;
		word[15'd1530] <= 32'd606;
		word[15'd1531] <= 32'd607;
		word[15'd1532] <= 32'd608;
		word[15'd1533] <= 32'd609;
		word[15'd1534] <= 32'd610;
		word[15'd1535] <= 32'd611;
		word[15'd1536] <= 32'd612;
		word[15'd1537] <= 32'd613;
		word[15'd1538] <= 32'd614;
		word[15'd1539] <= 32'd615;
		word[15'd1540] <= 32'd616;
		word[15'd1541] <= 32'd617;
		word[15'd1542] <= 32'd618;
		word[15'd1543] <= 32'd619;
		word[15'd1544] <= 32'd620;
		word[15'd1545] <= 32'd621;
		word[15'd1546] <= 32'd622;
		word[15'd1547] <= 32'd623;
		word[15'd1548] <= 32'd624;
		word[15'd1549] <= 32'd625;
		word[15'd1550] <= 32'd626;
		word[15'd1551] <= 32'd627;
		word[15'd1552] <= 32'd628;
		word[15'd1553] <= 32'd629;
		word[15'd1554] <= 32'd630;
		word[15'd1555] <= 32'd631;
		word[15'd1556] <= 32'd632;
		word[15'd1557] <= 32'd633;
		word[15'd1558] <= 32'd634;
		word[15'd1559] <= 32'd635;
		word[15'd1560] <= 32'd636;
		word[15'd1561] <= 32'd637;
		word[15'd1562] <= 32'd638;
		word[15'd1563] <= 32'd639;
		word[15'd1564] <= 32'd640;
		word[15'd1565] <= 32'd641;
		word[15'd1566] <= 32'd642;
		word[15'd1567] <= 32'd643;
		word[15'd1568] <= 32'd644;
		word[15'd1569] <= 32'd645;
		word[15'd1570] <= 32'd646;
		word[15'd1571] <= 32'd647;
		word[15'd1572] <= 32'd648;
		word[15'd1573] <= 32'd649;
		word[15'd1574] <= 32'd650;
		word[15'd1575] <= 32'd651;
		word[15'd1576] <= 32'd652;
		word[15'd1577] <= 32'd653;
		word[15'd1578] <= 32'd654;
		word[15'd1579] <= 32'd655;
		word[15'd1580] <= 32'd656;
		word[15'd1581] <= 32'd657;
		word[15'd1582] <= 32'd658;
		word[15'd1583] <= 32'd659;
		word[15'd1584] <= 32'd660;
		word[15'd1585] <= 32'd661;
		word[15'd1586] <= 32'd662;
		word[15'd1587] <= 32'd663;
		word[15'd1588] <= 32'd664;
		word[15'd1589] <= 32'd665;
		word[15'd1590] <= 32'd666;
		word[15'd1591] <= 32'd667;
		word[15'd1592] <= 32'd668;
		word[15'd1593] <= 32'd669;
		word[15'd1594] <= 32'd670;
		word[15'd1595] <= 32'd671;
		word[15'd1596] <= 32'd672;
		word[15'd1597] <= 32'd673;
		word[15'd1598] <= 32'd674;
		word[15'd1599] <= 32'd675;
		word[15'd1600] <= 32'd676;
		word[15'd1601] <= 32'd677;
		word[15'd1602] <= 32'd678;
		word[15'd1603] <= 32'd679;
		word[15'd1604] <= 32'd680;
		word[15'd1605] <= 32'd681;
		word[15'd1606] <= 32'd682;
		word[15'd1607] <= 32'd683;
		word[15'd1608] <= 32'd684;
		word[15'd1609] <= 32'd685;
		word[15'd1610] <= 32'd686;
		word[15'd1611] <= 32'd687;
		word[15'd1612] <= 32'd688;
		word[15'd1613] <= 32'd689;
		word[15'd1614] <= 32'd690;
		word[15'd1615] <= 32'd691;
		word[15'd1616] <= 32'd692;
		word[15'd1617] <= 32'd693;
		word[15'd1618] <= 32'd694;
		word[15'd1619] <= 32'd695;
		word[15'd1620] <= 32'd696;
		word[15'd1621] <= 32'd697;
		word[15'd1622] <= 32'd698;
		word[15'd1623] <= 32'd699;
		word[15'd1624] <= 32'd700;
		word[15'd1625] <= 32'd701;
		word[15'd1626] <= 32'd702;
		word[15'd1627] <= 32'd703;
		word[15'd1628] <= 32'd704;
		word[15'd1629] <= 32'd705;
		word[15'd1630] <= 32'd706;
		word[15'd1631] <= 32'd707;
		word[15'd1632] <= 32'd708;
		word[15'd1633] <= 32'd709;
		word[15'd1634] <= 32'd710;
		word[15'd1635] <= 32'd711;
		word[15'd1636] <= 32'd712;
		word[15'd1637] <= 32'd713;
		word[15'd1638] <= 32'd714;
		word[15'd1639] <= 32'd715;
		word[15'd1640] <= 32'd716;
		word[15'd1641] <= 32'd717;
		word[15'd1642] <= 32'd718;
		word[15'd1643] <= 32'd719;
		word[15'd1644] <= 32'd720;
		word[15'd1645] <= 32'd721;
		word[15'd1646] <= 32'd722;
		word[15'd1647] <= 32'd723;
		word[15'd1648] <= 32'd724;
		word[15'd1649] <= 32'd725;
		word[15'd1650] <= 32'd726;
		word[15'd1651] <= 32'd727;
		word[15'd1652] <= 32'd728;
		word[15'd1653] <= 32'd729;
		word[15'd1654] <= 32'd730;
		word[15'd1655] <= 32'd731;
		word[15'd1656] <= 32'd732;
		word[15'd1657] <= 32'd733;
		word[15'd1658] <= 32'd734;
		word[15'd1659] <= 32'd735;
		word[15'd1660] <= 32'd736;
		word[15'd1661] <= 32'd737;
		word[15'd1662] <= 32'd738;
		word[15'd1663] <= 32'd739;
		word[15'd1664] <= 32'd740;
		word[15'd1665] <= 32'd741;
		word[15'd1666] <= 32'd742;
		word[15'd1667] <= 32'd743;
		word[15'd1668] <= 32'd744;
		word[15'd1669] <= 32'd745;
		word[15'd1670] <= 32'd746;
		word[15'd1671] <= 32'd747;
		word[15'd1672] <= 32'd748;
		word[15'd1673] <= 32'd749;
		word[15'd1674] <= 32'd750;
		word[15'd1675] <= 32'd751;
		word[15'd1676] <= 32'd752;
		word[15'd1677] <= 32'd753;
		word[15'd1678] <= 32'd754;
		word[15'd1679] <= 32'd755;
		word[15'd1680] <= 32'd756;
		word[15'd1681] <= 32'd757;
		word[15'd1682] <= 32'd758;
		word[15'd1683] <= 32'd759;
		word[15'd1684] <= 32'd760;
		word[15'd1685] <= 32'd761;
		word[15'd1686] <= 32'd762;
		word[15'd1687] <= 32'd763;
		word[15'd1688] <= 32'd764;
		word[15'd1689] <= 32'd765;
		word[15'd1690] <= 32'd766;
		word[15'd1691] <= 32'd767;
		word[15'd1692] <= 32'd768;
		word[15'd1693] <= 32'd769;
		word[15'd1694] <= 32'd770;
		word[15'd1695] <= 32'd771;
		word[15'd1696] <= 32'd772;
		word[15'd1697] <= 32'd773;
		word[15'd1698] <= 32'd774;
		word[15'd1699] <= 32'd775;
		word[15'd1700] <= 32'd776;
		word[15'd1701] <= 32'd777;
		word[15'd1702] <= 32'd778;
		word[15'd1703] <= 32'd779;
		word[15'd1704] <= 32'd780;
		word[15'd1705] <= 32'd781;
		word[15'd1706] <= 32'd782;
		word[15'd1707] <= 32'd783;
		word[15'd1708] <= 32'd784;
		word[15'd1709] <= 32'd785;
		word[15'd1710] <= 32'd786;
		word[15'd1711] <= 32'd787;
		word[15'd1712] <= 32'd788;
		word[15'd1713] <= 32'd789;
		word[15'd1714] <= 32'd790;
		word[15'd1715] <= 32'd791;
		word[15'd1716] <= 32'd792;
		word[15'd1717] <= 32'd793;
		word[15'd1718] <= 32'd794;
		word[15'd1719] <= 32'd795;
		word[15'd1720] <= 32'd796;
		word[15'd1721] <= 32'd797;
		word[15'd1722] <= 32'd798;
		word[15'd1723] <= 32'd799;
		word[15'd1724] <= 32'd800;
		word[15'd1725] <= 32'd801;
		word[15'd1726] <= 32'd802;
		word[15'd1727] <= 32'd803;
		word[15'd1728] <= 32'd804;
		word[15'd1729] <= 32'd805;
		word[15'd1730] <= 32'd806;
		word[15'd1731] <= 32'd807;
		word[15'd1732] <= 32'd808;
		word[15'd1733] <= 32'd809;
		word[15'd1734] <= 32'd810;
		word[15'd1735] <= 32'd811;
		word[15'd1736] <= 32'd812;
		word[15'd1737] <= 32'd813;
		word[15'd1738] <= 32'd814;
		word[15'd1739] <= 32'd815;
		word[15'd1740] <= 32'd816;
		word[15'd1741] <= 32'd817;
		word[15'd1742] <= 32'd818;
		word[15'd1743] <= 32'd819;
		word[15'd1744] <= 32'd820;
		word[15'd1745] <= 32'd821;
		word[15'd1746] <= 32'd822;
		word[15'd1747] <= 32'd823;
		word[15'd1748] <= 32'd824;
		word[15'd1749] <= 32'd825;
		word[15'd1750] <= 32'd826;
		word[15'd1751] <= 32'd827;
		word[15'd1752] <= 32'd828;
		word[15'd1753] <= 32'd829;
		word[15'd1754] <= 32'd830;
		word[15'd1755] <= 32'd831;
		word[15'd1756] <= 32'd832;
		word[15'd1757] <= 32'd833;
		word[15'd1758] <= 32'd834;
		word[15'd1759] <= 32'd835;
		word[15'd1760] <= 32'd836;
		word[15'd1761] <= 32'd837;
		word[15'd1762] <= 32'd838;
		word[15'd1763] <= 32'd839;
		word[15'd1764] <= 32'd840;
		word[15'd1765] <= 32'd841;
		word[15'd1766] <= 32'd842;
		word[15'd1767] <= 32'd843;
		word[15'd1768] <= 32'd844;
		word[15'd1769] <= 32'd845;
		word[15'd1770] <= 32'd846;
		word[15'd1771] <= 32'd847;
		word[15'd1772] <= 32'd848;
		word[15'd1773] <= 32'd849;
		word[15'd1774] <= 32'd850;
		word[15'd1775] <= 32'd851;
		word[15'd1776] <= 32'd852;
		word[15'd1777] <= 32'd853;
		word[15'd1778] <= 32'd854;
		word[15'd1779] <= 32'd855;
		word[15'd1780] <= 32'd856;
		word[15'd1781] <= 32'd857;
		word[15'd1782] <= 32'd858;
		word[15'd1783] <= 32'd859;
		word[15'd1784] <= 32'd860;
		word[15'd1785] <= 32'd861;
		word[15'd1786] <= 32'd862;
		word[15'd1787] <= 32'd863;
		word[15'd1788] <= 32'd864;
		word[15'd1789] <= 32'd865;
		word[15'd1790] <= 32'd866;
		word[15'd1791] <= 32'd867;
		word[15'd1792] <= 32'd868;
		word[15'd1793] <= 32'd869;
		word[15'd1794] <= 32'd870;
		word[15'd1795] <= 32'd871;
		word[15'd1796] <= 32'd872;
		word[15'd1797] <= 32'd873;
		word[15'd1798] <= 32'd874;
		word[15'd1799] <= 32'd875;
		word[15'd1800] <= 32'd876;
		word[15'd1801] <= 32'd877;
		word[15'd1802] <= 32'd878;
		word[15'd1803] <= 32'd879;
		word[15'd1804] <= 32'd880;
		word[15'd1805] <= 32'd881;
		word[15'd1806] <= 32'd882;
		word[15'd1807] <= 32'd883;
		word[15'd1808] <= 32'd884;
		word[15'd1809] <= 32'd885;
		word[15'd1810] <= 32'd886;
		word[15'd1811] <= 32'd887;
		word[15'd1812] <= 32'd888;
		word[15'd1813] <= 32'd889;
		word[15'd1814] <= 32'd890;
		word[15'd1815] <= 32'd891;
		word[15'd1816] <= 32'd892;
		word[15'd1817] <= 32'd893;
		word[15'd1818] <= 32'd894;
		word[15'd1819] <= 32'd895;
		word[15'd1820] <= 32'd896;
		word[15'd1821] <= 32'd897;
		word[15'd1822] <= 32'd898;
		word[15'd1823] <= 32'd899;
		word[15'd1824] <= 32'd900;
		word[15'd1825] <= 32'd901;
		word[15'd1826] <= 32'd902;
		word[15'd1827] <= 32'd903;
		word[15'd1828] <= 32'd904;
		word[15'd1829] <= 32'd905;
		word[15'd1830] <= 32'd906;
		word[15'd1831] <= 32'd907;
		word[15'd1832] <= 32'd908;
		word[15'd1833] <= 32'd909;
		word[15'd1834] <= 32'd910;
		word[15'd1835] <= 32'd911;
		word[15'd1836] <= 32'd912;
		word[15'd1837] <= 32'd913;
		word[15'd1838] <= 32'd914;
		word[15'd1839] <= 32'd915;
		word[15'd1840] <= 32'd916;
		word[15'd1841] <= 32'd917;
		word[15'd1842] <= 32'd918;
		word[15'd1843] <= 32'd919;
		word[15'd1844] <= 32'd920;
		word[15'd1845] <= 32'd921;
		word[15'd1846] <= 32'd922;
		word[15'd1847] <= 32'd923;
		word[15'd1848] <= 32'd924;
		word[15'd1849] <= 32'd925;
		word[15'd1850] <= 32'd926;
		word[15'd1851] <= 32'd927;
		word[15'd1852] <= 32'd928;
		word[15'd1853] <= 32'd929;
		word[15'd1854] <= 32'd930;
		word[15'd1855] <= 32'd931;
		word[15'd1856] <= 32'd932;
		word[15'd1857] <= 32'd933;
		word[15'd1858] <= 32'd934;
		word[15'd1859] <= 32'd935;
		word[15'd1860] <= 32'd936;
		word[15'd1861] <= 32'd937;
		word[15'd1862] <= 32'd938;
		word[15'd1863] <= 32'd939;
		word[15'd1864] <= 32'd940;
		word[15'd1865] <= 32'd941;
		word[15'd1866] <= 32'd942;
		word[15'd1867] <= 32'd943;
		word[15'd1868] <= 32'd944;
		word[15'd1869] <= 32'd945;
		word[15'd1870] <= 32'd946;
		word[15'd1871] <= 32'd947;
		word[15'd1872] <= 32'd948;
		word[15'd1873] <= 32'd949;
		word[15'd1874] <= 32'd950;
		word[15'd1875] <= 32'd951;
		word[15'd1876] <= 32'd952;
		word[15'd1877] <= 32'd953;
		word[15'd1878] <= 32'd954;
		word[15'd1879] <= 32'd955;
		word[15'd1880] <= 32'd956;
		word[15'd1881] <= 32'd957;
		word[15'd1882] <= 32'd958;
		word[15'd1883] <= 32'd959;
		word[15'd1884] <= 32'd960;
		word[15'd1885] <= 32'd961;
		word[15'd1886] <= 32'd962;
		word[15'd1887] <= 32'd963;
		word[15'd1888] <= 32'd964;
		word[15'd1889] <= 32'd965;
		word[15'd1890] <= 32'd966;
		word[15'd1891] <= 32'd967;
		word[15'd1892] <= 32'd968;
		word[15'd1893] <= 32'd969;
		word[15'd1894] <= 32'd970;
		word[15'd1895] <= 32'd971;
		word[15'd1896] <= 32'd972;
		word[15'd1897] <= 32'd973;
		word[15'd1898] <= 32'd974;
		word[15'd1899] <= 32'd975;
		word[15'd1900] <= 32'd976;
		word[15'd1901] <= 32'd977;
		word[15'd1902] <= 32'd978;
		word[15'd1903] <= 32'd979;
		word[15'd1904] <= 32'd980;
		word[15'd1905] <= 32'd981;
		word[15'd1906] <= 32'd982;
		word[15'd1907] <= 32'd983;
		word[15'd1908] <= 32'd984;
		word[15'd1909] <= 32'd985;
		word[15'd1910] <= 32'd986;
		word[15'd1911] <= 32'd987;
		word[15'd1912] <= 32'd988;
		word[15'd1913] <= 32'd989;
		word[15'd1914] <= 32'd990;
		word[15'd1915] <= 32'd991;
		word[15'd1916] <= 32'd992;
		word[15'd1917] <= 32'd993;
		word[15'd1918] <= 32'd994;
		word[15'd1919] <= 32'd995;
		word[15'd1920] <= 32'd996;
		word[15'd1921] <= 32'd997;
		word[15'd1922] <= 32'd998;
		word[15'd1923] <= 32'd999;
		word[15'd1924] <= 32'd1000;
		word[15'd1925] <= 32'd1001;
		word[15'd1926] <= 32'd1002;
		word[15'd1927] <= 32'd1003;
		word[15'd1928] <= 32'd1004;
		word[15'd1929] <= 32'd1005;
		word[15'd1930] <= 32'd1006;
		word[15'd1931] <= 32'd1007;
		word[15'd1932] <= 32'd1008;
		word[15'd1933] <= 32'd1009;
		word[15'd1934] <= 32'd1010;
		word[15'd1935] <= 32'd1011;
		word[15'd1936] <= 32'd1012;
		word[15'd1937] <= 32'd1013;
		word[15'd1938] <= 32'd1014;
		word[15'd1939] <= 32'd1015;
		word[15'd1940] <= 32'd1016;
		word[15'd1941] <= 32'd1017;
		word[15'd1942] <= 32'd1018;
		word[15'd1943] <= 32'd1019;
		word[15'd1944] <= 32'd1020;
		word[15'd1945] <= 32'd1021;
		word[15'd1946] <= 32'd1022;
		word[15'd1947] <= 32'd1023;
		word[15'd1948] <= 32'd1024;
		word[15'd1949] <= 32'd1025;
		word[15'd1950] <= 32'd1026;
		word[15'd1951] <= 32'd1027;
		word[15'd1952] <= 32'd1028;
		word[15'd1953] <= 32'd1029;
		word[15'd1954] <= 32'd1030;
		word[15'd1955] <= 32'd1031;
		word[15'd1956] <= 32'd1032;
		word[15'd1957] <= 32'd1033;
		word[15'd1958] <= 32'd1034;
		word[15'd1959] <= 32'd1035;
		word[15'd1960] <= 32'd1036;
		word[15'd1961] <= 32'd1037;
		word[15'd1962] <= 32'd1038;
		word[15'd1963] <= 32'd1039;
		word[15'd1964] <= 32'd1040;
		word[15'd1965] <= 32'd1041;
		word[15'd1966] <= 32'd1042;
		word[15'd1967] <= 32'd1043;
		word[15'd1968] <= 32'd1044;
		word[15'd1969] <= 32'd1045;
		word[15'd1970] <= 32'd1046;
		word[15'd1971] <= 32'd1047;
		word[15'd1972] <= 32'd1048;
		word[15'd1973] <= 32'd1049;
		word[15'd1974] <= 32'd1050;
		word[15'd1975] <= 32'd1051;
		word[15'd1976] <= 32'd1052;
		word[15'd1977] <= 32'd1053;
		word[15'd1978] <= 32'd1054;
		word[15'd1979] <= 32'd1055;
		word[15'd1980] <= 32'd1056;
		word[15'd1981] <= 32'd1057;
		word[15'd1982] <= 32'd1058;
		word[15'd1983] <= 32'd1059;
		word[15'd1984] <= 32'd1060;
		word[15'd1985] <= 32'd1061;
		word[15'd1986] <= 32'd1062;
		word[15'd1987] <= 32'd1063;
		word[15'd1988] <= 32'd1064;
		word[15'd1989] <= 32'd1065;
		word[15'd1990] <= 32'd1066;
		word[15'd1991] <= 32'd1067;
		word[15'd1992] <= 32'd1068;
		word[15'd1993] <= 32'd1069;
		word[15'd1994] <= 32'd1070;
		word[15'd1995] <= 32'd1071;
		word[15'd1996] <= 32'd1072;
		word[15'd1997] <= 32'd1073;
		word[15'd1998] <= 32'd1074;
		word[15'd1999] <= 32'd1075;
		word[15'd2000] <= 32'd1076;
		word[15'd2001] <= 32'd1077;
		word[15'd2002] <= 32'd1078;
		word[15'd2003] <= 32'd1079;
		word[15'd2004] <= 32'd1080;
		word[15'd2005] <= 32'd1081;
		word[15'd2006] <= 32'd1082;
		word[15'd2007] <= 32'd1083;
		word[15'd2008] <= 32'd1084;
		word[15'd2009] <= 32'd1085;
		word[15'd2010] <= 32'd1086;
		word[15'd2011] <= 32'd1087;
		word[15'd2012] <= 32'd1088;
		word[15'd2013] <= 32'd1089;
		word[15'd2014] <= 32'd1090;
		word[15'd2015] <= 32'd1091;
		word[15'd2016] <= 32'd1092;
		word[15'd2017] <= 32'd1093;
		word[15'd2018] <= 32'd1094;
		word[15'd2019] <= 32'd1095;
		word[15'd2020] <= 32'd1096;
		word[15'd2021] <= 32'd1097;
		word[15'd2022] <= 32'd1098;
		word[15'd2023] <= 32'd1099;
		word[15'd2024] <= 32'd1100;
		word[15'd2025] <= 32'd1101;
		word[15'd2026] <= 32'd1102;
		word[15'd2027] <= 32'd1103;
		word[15'd2028] <= 32'd1104;
		word[15'd2029] <= 32'd1105;
		word[15'd2030] <= 32'd1106;
		word[15'd2031] <= 32'd1107;
		word[15'd2032] <= 32'd1108;
		word[15'd2033] <= 32'd1109;
		word[15'd2034] <= 32'd1110;
		word[15'd2035] <= 32'd1111;
		word[15'd2036] <= 32'd1112;
		word[15'd2037] <= 32'd1113;
		word[15'd2038] <= 32'd1114;
		word[15'd2039] <= 32'd1115;
		word[15'd2040] <= 32'd1116;
		word[15'd2041] <= 32'd1117;
		word[15'd2042] <= 32'd1118;
		word[15'd2043] <= 32'd1119;
		word[15'd2044] <= 32'd1120;
		word[15'd2045] <= 32'd1121;
		word[15'd2046] <= 32'd1122;
		word[15'd2047] <= 32'd1123;
		word[15'd2048] <= 32'd1124;
		word[15'd2049] <= 32'd1125;
		word[15'd2050] <= 32'd1126;
		word[15'd2051] <= 32'd1127;
		word[15'd2052] <= 32'd1128;
		word[15'd2053] <= 32'd1129;
		word[15'd2054] <= 32'd1130;
		word[15'd2055] <= 32'd1131;
		word[15'd2056] <= 32'd1132;
		word[15'd2057] <= 32'd1133;
		word[15'd2058] <= 32'd1134;
		word[15'd2059] <= 32'd1135;
		word[15'd2060] <= 32'd1136;
		word[15'd2061] <= 32'd1137;
		word[15'd2062] <= 32'd1138;
		word[15'd2063] <= 32'd1139;
		word[15'd2064] <= 32'd1140;
		word[15'd2065] <= 32'd1141;
		word[15'd2066] <= 32'd1142;
		word[15'd2067] <= 32'd1143;
		word[15'd2068] <= 32'd1144;
		word[15'd2069] <= 32'd1145;
		word[15'd2070] <= 32'd1146;
		word[15'd2071] <= 32'd1147;
		word[15'd2072] <= 32'd1148;
		word[15'd2073] <= 32'd1149;
		word[15'd2074] <= 32'd1150;
		word[15'd2075] <= 32'd1151;
		word[15'd2076] <= 32'd1152;
		word[15'd2077] <= 32'd1153;
		word[15'd2078] <= 32'd1154;
		word[15'd2079] <= 32'd1155;
		word[15'd2080] <= 32'd1156;
		word[15'd2081] <= 32'd1157;
		word[15'd2082] <= 32'd1158;
		word[15'd2083] <= 32'd1159;
		word[15'd2084] <= 32'd1160;
		word[15'd2085] <= 32'd1161;
		word[15'd2086] <= 32'd1162;
		word[15'd2087] <= 32'd1163;
		word[15'd2088] <= 32'd1164;
		word[15'd2089] <= 32'd1165;
		word[15'd2090] <= 32'd1166;
		word[15'd2091] <= 32'd1167;
		word[15'd2092] <= 32'd1168;
		word[15'd2093] <= 32'd1169;
		word[15'd2094] <= 32'd1170;
		word[15'd2095] <= 32'd1171;
		word[15'd2096] <= 32'd1172;
		word[15'd2097] <= 32'd1173;
		word[15'd2098] <= 32'd1174;
		word[15'd2099] <= 32'd1175;
		word[15'd2100] <= 32'd1176;
		word[15'd2101] <= 32'd1177;
		word[15'd2102] <= 32'd1178;
		word[15'd2103] <= 32'd1179;
		word[15'd2104] <= 32'd1180;
		word[15'd2105] <= 32'd1181;
		word[15'd2106] <= 32'd1182;
		word[15'd2107] <= 32'd1183;
		word[15'd2108] <= 32'd1184;
		word[15'd2109] <= 32'd1185;
		word[15'd2110] <= 32'd1186;
		word[15'd2111] <= 32'd1187;
		word[15'd2112] <= 32'd1188;
		word[15'd2113] <= 32'd1189;
		word[15'd2114] <= 32'd1190;
		word[15'd2115] <= 32'd1191;
		word[15'd2116] <= 32'd1192;
		word[15'd2117] <= 32'd1193;
		word[15'd2118] <= 32'd1194;
		word[15'd2119] <= 32'd1195;
		word[15'd2120] <= 32'd1196;
		word[15'd2121] <= 32'd1197;
		word[15'd2122] <= 32'd1198;
		word[15'd2123] <= 32'd1199;
		word[15'd2124] <= 32'd1200;
		word[15'd2125] <= 32'd1201;
		word[15'd2126] <= 32'd1202;
		word[15'd2127] <= 32'd1203;
		word[15'd2128] <= 32'd1204;
		word[15'd2129] <= 32'd1205;
		word[15'd2130] <= 32'd1206;
		word[15'd2131] <= 32'd1207;
		word[15'd2132] <= 32'd1208;
		word[15'd2133] <= 32'd1209;
		word[15'd2134] <= 32'd1210;
		word[15'd2135] <= 32'd1211;
		word[15'd2136] <= 32'd1212;
		word[15'd2137] <= 32'd1213;
		word[15'd2138] <= 32'd1214;
		word[15'd2139] <= 32'd1215;
		word[15'd2140] <= 32'd1216;
		word[15'd2141] <= 32'd1217;
		word[15'd2142] <= 32'd1218;
		word[15'd2143] <= 32'd1219;
		word[15'd2144] <= 32'd1220;
		word[15'd2145] <= 32'd1221;
		word[15'd2146] <= 32'd1222;
		word[15'd2147] <= 32'd1223;
		word[15'd2148] <= 32'd1224;
		word[15'd2149] <= 32'd1225;
		word[15'd2150] <= 32'd1226;
		word[15'd2151] <= 32'd1227;
		word[15'd2152] <= 32'd1228;
		word[15'd2153] <= 32'd1229;
		word[15'd2154] <= 32'd1230;
		word[15'd2155] <= 32'd1231;
		word[15'd2156] <= 32'd1232;
		word[15'd2157] <= 32'd1233;
		word[15'd2158] <= 32'd1234;
		word[15'd2159] <= 32'd1235;
		word[15'd2160] <= 32'd1236;
		word[15'd2161] <= 32'd1237;
		word[15'd2162] <= 32'd1238;
		word[15'd2163] <= 32'd1239;
		word[15'd2164] <= 32'd1240;
		word[15'd2165] <= 32'd1241;
		word[15'd2166] <= 32'd1242;
		word[15'd2167] <= 32'd1243;
		word[15'd2168] <= 32'd1244;
		word[15'd2169] <= 32'd1245;
		word[15'd2170] <= 32'd1246;
		word[15'd2171] <= 32'd1247;
		word[15'd2172] <= 32'd1248;
		word[15'd2173] <= 32'd1249;
		word[15'd2174] <= 32'd1250;
		word[15'd2175] <= 32'd1251;
		word[15'd2176] <= 32'd1252;
		word[15'd2177] <= 32'd1253;
		word[15'd2178] <= 32'd1254;
		word[15'd2179] <= 32'd1255;
		word[15'd2180] <= 32'd1256;
		word[15'd2181] <= 32'd1257;
		word[15'd2182] <= 32'd1258;
		word[15'd2183] <= 32'd1259;
		word[15'd2184] <= 32'd1260;
		word[15'd2185] <= 32'd1261;
		word[15'd2186] <= 32'd1262;
		word[15'd2187] <= 32'd1263;
		word[15'd2188] <= 32'd1264;
		word[15'd2189] <= 32'd1265;
		word[15'd2190] <= 32'd1266;
		word[15'd2191] <= 32'd1267;
		word[15'd2192] <= 32'd1268;
		word[15'd2193] <= 32'd1269;
		word[15'd2194] <= 32'd1270;
		word[15'd2195] <= 32'd1271;
		word[15'd2196] <= 32'd1272;
		word[15'd2197] <= 32'd1273;
		word[15'd2198] <= 32'd1274;
		word[15'd2199] <= 32'd1275;
		word[15'd2200] <= 32'd1276;
		word[15'd2201] <= 32'd1277;
		word[15'd2202] <= 32'd1278;
		word[15'd2203] <= 32'd1279;
		word[15'd2204] <= 32'd1280;
		word[15'd2205] <= 32'd1281;
		word[15'd2206] <= 32'd1282;
		word[15'd2207] <= 32'd1283;
		word[15'd2208] <= 32'd1284;
		word[15'd2209] <= 32'd1285;
		word[15'd2210] <= 32'd1286;
		word[15'd2211] <= 32'd1287;
		word[15'd2212] <= 32'd1288;
		word[15'd2213] <= 32'd1289;
		word[15'd2214] <= 32'd1290;
		word[15'd2215] <= 32'd1291;
		word[15'd2216] <= 32'd1292;
		word[15'd2217] <= 32'd1293;
		word[15'd2218] <= 32'd1294;
		word[15'd2219] <= 32'd1295;
		word[15'd2220] <= 32'd1296;
		word[15'd2221] <= 32'd1297;
		word[15'd2222] <= 32'd1298;
		word[15'd2223] <= 32'd1299;
		word[15'd2224] <= 32'd1300;
		word[15'd2225] <= 32'd1301;
		word[15'd2226] <= 32'd1302;
		word[15'd2227] <= 32'd1303;
		word[15'd2228] <= 32'd1304;
		word[15'd2229] <= 32'd1305;
		word[15'd2230] <= 32'd1306;
		word[15'd2231] <= 32'd1307;
		word[15'd2232] <= 32'd1308;
		word[15'd2233] <= 32'd1309;
		word[15'd2234] <= 32'd1310;
		word[15'd2235] <= 32'd1311;
		word[15'd2236] <= 32'd1312;
		word[15'd2237] <= 32'd1313;
		word[15'd2238] <= 32'd1314;
		word[15'd2239] <= 32'd1315;
		word[15'd2240] <= 32'd1316;
		word[15'd2241] <= 32'd1317;
		word[15'd2242] <= 32'd1318;
		word[15'd2243] <= 32'd1319;
		word[15'd2244] <= 32'd1320;
		word[15'd2245] <= 32'd1321;
		word[15'd2246] <= 32'd1322;
		word[15'd2247] <= 32'd1323;
		word[15'd2248] <= 32'd1324;
		word[15'd2249] <= 32'd1325;
		word[15'd2250] <= 32'd1326;
		word[15'd2251] <= 32'd1327;
		word[15'd2252] <= 32'd1328;
		word[15'd2253] <= 32'd1329;
		word[15'd2254] <= 32'd1330;
		word[15'd2255] <= 32'd1331;
		word[15'd2256] <= 32'd1332;
		word[15'd2257] <= 32'd1333;
		word[15'd2258] <= 32'd1334;
		word[15'd2259] <= 32'd1335;
		word[15'd2260] <= 32'd1336;
		word[15'd2261] <= 32'd1337;
		word[15'd2262] <= 32'd1338;
		word[15'd2263] <= 32'd1339;
		word[15'd2264] <= 32'd1340;
		word[15'd2265] <= 32'd1341;
		word[15'd2266] <= 32'd1342;
		word[15'd2267] <= 32'd1343;
		word[15'd2268] <= 32'd1344;
		word[15'd2269] <= 32'd1345;
		word[15'd2270] <= 32'd1346;
		word[15'd2271] <= 32'd1347;
		word[15'd2272] <= 32'd1348;
		word[15'd2273] <= 32'd1349;
		word[15'd2274] <= 32'd1350;
		word[15'd2275] <= 32'd1351;
		word[15'd2276] <= 32'd1352;
		word[15'd2277] <= 32'd1353;
		word[15'd2278] <= 32'd1354;
		word[15'd2279] <= 32'd1355;
		word[15'd2280] <= 32'd1356;
		word[15'd2281] <= 32'd1357;
		word[15'd2282] <= 32'd1358;
		word[15'd2283] <= 32'd1359;
		word[15'd2284] <= 32'd1360;
		word[15'd2285] <= 32'd1361;
		word[15'd2286] <= 32'd1362;
		word[15'd2287] <= 32'd1363;
		word[15'd2288] <= 32'd1364;
		word[15'd2289] <= 32'd1365;
		word[15'd2290] <= 32'd1366;
		word[15'd2291] <= 32'd1367;
		word[15'd2292] <= 32'd1368;
		word[15'd2293] <= 32'd1369;
		word[15'd2294] <= 32'd1370;
		word[15'd2295] <= 32'd1371;
		word[15'd2296] <= 32'd1372;
		word[15'd2297] <= 32'd1373;
		word[15'd2298] <= 32'd1374;
		word[15'd2299] <= 32'd1375;
		word[15'd2300] <= 32'd1376;
		word[15'd2301] <= 32'd1377;
		word[15'd2302] <= 32'd1378;
		word[15'd2303] <= 32'd1379;
		word[15'd2304] <= 32'd1380;
		word[15'd2305] <= 32'd1381;
		word[15'd2306] <= 32'd1382;
		word[15'd2307] <= 32'd1383;
		word[15'd2308] <= 32'd1384;
		word[15'd2309] <= 32'd1385;
		word[15'd2310] <= 32'd1386;
		word[15'd2311] <= 32'd1387;
		word[15'd2312] <= 32'd1388;
		word[15'd2313] <= 32'd1389;
		word[15'd2314] <= 32'd1390;
		word[15'd2315] <= 32'd1391;
		word[15'd2316] <= 32'd1392;
		word[15'd2317] <= 32'd1393;
		word[15'd2318] <= 32'd1394;
		word[15'd2319] <= 32'd1395;
		word[15'd2320] <= 32'd1396;
		word[15'd2321] <= 32'd1397;
		word[15'd2322] <= 32'd1398;
		word[15'd2323] <= 32'd1399;
		word[15'd2324] <= 32'd1400;
		word[15'd2325] <= 32'd1401;
		word[15'd2326] <= 32'd1402;
		word[15'd2327] <= 32'd1403;
		word[15'd2328] <= 32'd1404;
		word[15'd2329] <= 32'd1405;
		word[15'd2330] <= 32'd1406;
		word[15'd2331] <= 32'd1407;
		word[15'd2332] <= 32'd1408;
		word[15'd2333] <= 32'd1409;
		word[15'd2334] <= 32'd1410;
		word[15'd2335] <= 32'd1411;
		word[15'd2336] <= 32'd1412;
		word[15'd2337] <= 32'd1413;
		word[15'd2338] <= 32'd1414;
		word[15'd2339] <= 32'd1415;
		word[15'd2340] <= 32'd1416;
		word[15'd2341] <= 32'd1417;
		word[15'd2342] <= 32'd1418;
		word[15'd2343] <= 32'd1419;
		word[15'd2344] <= 32'd1420;
		word[15'd2345] <= 32'd1421;
		word[15'd2346] <= 32'd1422;
		word[15'd2347] <= 32'd1423;
		word[15'd2348] <= 32'd1424;
		word[15'd2349] <= 32'd1425;
		word[15'd2350] <= 32'd1426;
		word[15'd2351] <= 32'd1427;
		word[15'd2352] <= 32'd1428;
		word[15'd2353] <= 32'd1429;
		word[15'd2354] <= 32'd1430;
		word[15'd2355] <= 32'd1431;
		word[15'd2356] <= 32'd1432;
		word[15'd2357] <= 32'd1433;
		word[15'd2358] <= 32'd1434;
		word[15'd2359] <= 32'd1435;
		word[15'd2360] <= 32'd1436;
		word[15'd2361] <= 32'd1437;
		word[15'd2362] <= 32'd1438;
		word[15'd2363] <= 32'd1439;
		word[15'd2364] <= 32'd1440;
		word[15'd2365] <= 32'd1441;
		word[15'd2366] <= 32'd1442;
		word[15'd2367] <= 32'd1443;
		word[15'd2368] <= 32'd1444;
		word[15'd2369] <= 32'd1445;
		word[15'd2370] <= 32'd1446;
		word[15'd2371] <= 32'd1447;
		word[15'd2372] <= 32'd1448;
		word[15'd2373] <= 32'd1449;
		word[15'd2374] <= 32'd1450;
		word[15'd2375] <= 32'd1451;
		word[15'd2376] <= 32'd1452;
		word[15'd2377] <= 32'd1453;
		word[15'd2378] <= 32'd1454;
		word[15'd2379] <= 32'd1455;
		word[15'd2380] <= 32'd1456;
		word[15'd2381] <= 32'd1457;
		word[15'd2382] <= 32'd1458;
		word[15'd2383] <= 32'd1459;
		word[15'd2384] <= 32'd1460;
		word[15'd2385] <= 32'd1461;
		word[15'd2386] <= 32'd1462;
		word[15'd2387] <= 32'd1463;
		word[15'd2388] <= 32'd1464;
		word[15'd2389] <= 32'd1465;
		word[15'd2390] <= 32'd1466;
		word[15'd2391] <= 32'd1467;
		word[15'd2392] <= 32'd1468;
		word[15'd2393] <= 32'd1469;
		word[15'd2394] <= 32'd1470;
		word[15'd2395] <= 32'd1471;
		word[15'd2396] <= 32'd1472;
		word[15'd2397] <= 32'd1473;
		word[15'd2398] <= 32'd1474;
		word[15'd2399] <= 32'd1475;
		word[15'd2400] <= 32'd1476;
		word[15'd2401] <= 32'd1477;
		word[15'd2402] <= 32'd1478;
		word[15'd2403] <= 32'd1479;
		word[15'd2404] <= 32'd1480;
		word[15'd2405] <= 32'd1481;
		word[15'd2406] <= 32'd1482;
		word[15'd2407] <= 32'd1483;
		word[15'd2408] <= 32'd1484;
		word[15'd2409] <= 32'd1485;
		word[15'd2410] <= 32'd1486;
		word[15'd2411] <= 32'd1487;
		word[15'd2412] <= 32'd1488;
		word[15'd2413] <= 32'd1489;
		word[15'd2414] <= 32'd1490;
		word[15'd2415] <= 32'd1491;
		word[15'd2416] <= 32'd1492;
		word[15'd2417] <= 32'd1493;
		word[15'd2418] <= 32'd1494;
		word[15'd2419] <= 32'd1495;
		word[15'd2420] <= 32'd1496;
		word[15'd2421] <= 32'd1497;
		word[15'd2422] <= 32'd1498;
		word[15'd2423] <= 32'd1499;
		word[15'd2424] <= 32'd1500;
		word[15'd2425] <= 32'd1501;
		word[15'd2426] <= 32'd1502;
		word[15'd2427] <= 32'd1503;
		word[15'd2428] <= 32'd1504;
		word[15'd2429] <= 32'd1505;
		word[15'd2430] <= 32'd1506;
		word[15'd2431] <= 32'd1507;
		word[15'd2432] <= 32'd1508;
		word[15'd2433] <= 32'd1509;
		word[15'd2434] <= 32'd1510;
		word[15'd2435] <= 32'd1511;
		word[15'd2436] <= 32'd1512;
		word[15'd2437] <= 32'd1513;
		word[15'd2438] <= 32'd1514;
		word[15'd2439] <= 32'd1515;
		word[15'd2440] <= 32'd1516;
		word[15'd2441] <= 32'd1517;
		word[15'd2442] <= 32'd1518;
		word[15'd2443] <= 32'd1519;
		word[15'd2444] <= 32'd1520;
		word[15'd2445] <= 32'd1521;
		word[15'd2446] <= 32'd1522;
		word[15'd2447] <= 32'd1523;
		word[15'd2448] <= 32'd1524;
		word[15'd2449] <= 32'd1525;
		word[15'd2450] <= 32'd1526;
		word[15'd2451] <= 32'd1527;
		word[15'd2452] <= 32'd1528;
		word[15'd2453] <= 32'd1529;
		word[15'd2454] <= 32'd1530;
		word[15'd2455] <= 32'd1531;
		word[15'd2456] <= 32'd1532;
		word[15'd2457] <= 32'd1533;
		word[15'd2458] <= 32'd1534;
		word[15'd2459] <= 32'd1535;
		word[15'd2460] <= 32'd1536;
		word[15'd2461] <= 32'd1537;
		word[15'd2462] <= 32'd1538;
		word[15'd2463] <= 32'd1539;
		word[15'd2464] <= 32'd1540;
		word[15'd2465] <= 32'd1541;
		word[15'd2466] <= 32'd1542;
		word[15'd2467] <= 32'd1543;
		word[15'd2468] <= 32'd1544;
		word[15'd2469] <= 32'd1545;
		word[15'd2470] <= 32'd1546;
		word[15'd2471] <= 32'd1547;
		word[15'd2472] <= 32'd1548;
		word[15'd2473] <= 32'd1549;
		word[15'd2474] <= 32'd1550;
		word[15'd2475] <= 32'd1551;
		word[15'd2476] <= 32'd1552;
		word[15'd2477] <= 32'd1553;
		word[15'd2478] <= 32'd1554;
		word[15'd2479] <= 32'd1555;
		word[15'd2480] <= 32'd1556;
		word[15'd2481] <= 32'd1557;
		word[15'd2482] <= 32'd1558;
		word[15'd2483] <= 32'd1559;
		word[15'd2484] <= 32'd1560;
		word[15'd2485] <= 32'd1561;
		word[15'd2486] <= 32'd1562;
		word[15'd2487] <= 32'd1563;
		word[15'd2488] <= 32'd1564;
		word[15'd2489] <= 32'd1565;
		word[15'd2490] <= 32'd1566;
		word[15'd2491] <= 32'd1567;
		word[15'd2492] <= 32'd1568;
		word[15'd2493] <= 32'd1569;
		word[15'd2494] <= 32'd1570;
		word[15'd2495] <= 32'd1571;
		word[15'd2496] <= 32'd1572;
		word[15'd2497] <= 32'd1573;
		word[15'd2498] <= 32'd1574;
		word[15'd2499] <= 32'd1575;
		word[15'd2500] <= 32'd1576;
		word[15'd2501] <= 32'd1577;
		word[15'd2502] <= 32'd1578;
		word[15'd2503] <= 32'd1579;
		word[15'd2504] <= 32'd1580;
		word[15'd2505] <= 32'd1581;
		word[15'd2506] <= 32'd1582;
		word[15'd2507] <= 32'd1583;
		word[15'd2508] <= 32'd1584;
		word[15'd2509] <= 32'd1585;
		word[15'd2510] <= 32'd1586;
		word[15'd2511] <= 32'd1587;
		word[15'd2512] <= 32'd1588;
		word[15'd2513] <= 32'd1589;
		word[15'd2514] <= 32'd1590;
		word[15'd2515] <= 32'd1591;
		word[15'd2516] <= 32'd1592;
		word[15'd2517] <= 32'd1593;
		word[15'd2518] <= 32'd1594;
		word[15'd2519] <= 32'd1595;
		word[15'd2520] <= 32'd1596;
		word[15'd2521] <= 32'd1597;
		word[15'd2522] <= 32'd1598;
		word[15'd2523] <= 32'd1599;
		word[15'd2524] <= 32'd1600;
		word[15'd2525] <= 32'd1601;
		word[15'd2526] <= 32'd1602;
		word[15'd2527] <= 32'd1603;
		word[15'd2528] <= 32'd1604;
		word[15'd2529] <= 32'd1605;
		word[15'd2530] <= 32'd1606;
		word[15'd2531] <= 32'd1607;
		word[15'd2532] <= 32'd1608;
		word[15'd2533] <= 32'd1609;
		word[15'd2534] <= 32'd1610;
		word[15'd2535] <= 32'd1611;
		word[15'd2536] <= 32'd1612;
		word[15'd2537] <= 32'd1613;
		word[15'd2538] <= 32'd1614;
		word[15'd2539] <= 32'd1615;
		word[15'd2540] <= 32'd1616;
		word[15'd2541] <= 32'd1617;
		word[15'd2542] <= 32'd1618;
		word[15'd2543] <= 32'd1619;
		word[15'd2544] <= 32'd1620;
		word[15'd2545] <= 32'd1621;
		word[15'd2546] <= 32'd1622;
		word[15'd2547] <= 32'd1623;
		word[15'd2548] <= 32'd1624;
		word[15'd2549] <= 32'd1625;
		word[15'd2550] <= 32'd1626;
		word[15'd2551] <= 32'd1627;
		word[15'd2552] <= 32'd1628;
		word[15'd2553] <= 32'd1629;
		word[15'd2554] <= 32'd1630;
		word[15'd2555] <= 32'd1631;
		word[15'd2556] <= 32'd1632;
		word[15'd2557] <= 32'd1633;
		word[15'd2558] <= 32'd1634;
		word[15'd2559] <= 32'd1635;
		word[15'd2560] <= 32'd1636;
		word[15'd2561] <= 32'd1637;
		word[15'd2562] <= 32'd1638;
		word[15'd2563] <= 32'd1639;
		word[15'd2564] <= 32'd1640;
		word[15'd2565] <= 32'd1641;
		word[15'd2566] <= 32'd1642;
		word[15'd2567] <= 32'd1643;
		word[15'd2568] <= 32'd1644;
		word[15'd2569] <= 32'd1645;
		word[15'd2570] <= 32'd1646;
		word[15'd2571] <= 32'd1647;
		word[15'd2572] <= 32'd1648;
		word[15'd2573] <= 32'd1649;
		word[15'd2574] <= 32'd1650;
		word[15'd2575] <= 32'd1651;
		word[15'd2576] <= 32'd1652;
		word[15'd2577] <= 32'd1653;
		word[15'd2578] <= 32'd1654;
		word[15'd2579] <= 32'd1655;
		word[15'd2580] <= 32'd1656;
		word[15'd2581] <= 32'd1657;
		word[15'd2582] <= 32'd1658;
		word[15'd2583] <= 32'd1659;
		word[15'd2584] <= 32'd1660;
		word[15'd2585] <= 32'd1661;
		word[15'd2586] <= 32'd1662;
		word[15'd2587] <= 32'd1663;
		word[15'd2588] <= 32'd1664;
		word[15'd2589] <= 32'd1665;
		word[15'd2590] <= 32'd1666;
		word[15'd2591] <= 32'd1667;
		word[15'd2592] <= 32'd1668;
		word[15'd2593] <= 32'd1669;
		word[15'd2594] <= 32'd1670;
		word[15'd2595] <= 32'd1671;
		word[15'd2596] <= 32'd1672;
		word[15'd2597] <= 32'd1673;
		word[15'd2598] <= 32'd1674;
		word[15'd2599] <= 32'd1675;
		word[15'd2600] <= 32'd1676;
		word[15'd2601] <= 32'd1677;
		word[15'd2602] <= 32'd1678;
		word[15'd2603] <= 32'd1679;
		word[15'd2604] <= 32'd1680;
		word[15'd2605] <= 32'd1681;
		word[15'd2606] <= 32'd1682;
		word[15'd2607] <= 32'd1683;
		word[15'd2608] <= 32'd1684;
		word[15'd2609] <= 32'd1685;
		word[15'd2610] <= 32'd1686;
		word[15'd2611] <= 32'd1687;
		word[15'd2612] <= 32'd1688;
		word[15'd2613] <= 32'd1689;
		word[15'd2614] <= 32'd1690;
		word[15'd2615] <= 32'd1691;
		word[15'd2616] <= 32'd1692;
		word[15'd2617] <= 32'd1693;
		word[15'd2618] <= 32'd1694;
		word[15'd2619] <= 32'd1695;
		word[15'd2620] <= 32'd1696;
		word[15'd2621] <= 32'd1697;
		word[15'd2622] <= 32'd1698;
		word[15'd2623] <= 32'd1699;
		word[15'd2624] <= 32'd1700;
		word[15'd2625] <= 32'd1701;
		word[15'd2626] <= 32'd1702;
		word[15'd2627] <= 32'd1703;
		word[15'd2628] <= 32'd1704;
		word[15'd2629] <= 32'd1705;
		word[15'd2630] <= 32'd1706;
		word[15'd2631] <= 32'd1707;
		word[15'd2632] <= 32'd1708;
		word[15'd2633] <= 32'd1709;
		word[15'd2634] <= 32'd1710;
		word[15'd2635] <= 32'd1711;
		word[15'd2636] <= 32'd1712;
		word[15'd2637] <= 32'd1713;
		word[15'd2638] <= 32'd1714;
		word[15'd2639] <= 32'd1715;
		word[15'd2640] <= 32'd1716;
		word[15'd2641] <= 32'd1717;
		word[15'd2642] <= 32'd1718;
		word[15'd2643] <= 32'd1719;
		word[15'd2644] <= 32'd1720;
		word[15'd2645] <= 32'd1721;
		word[15'd2646] <= 32'd1722;
		word[15'd2647] <= 32'd1723;
		word[15'd2648] <= 32'd1724;
		word[15'd2649] <= 32'd1725;
		word[15'd2650] <= 32'd1726;
		word[15'd2651] <= 32'd1727;
		word[15'd2652] <= 32'd1728;
		word[15'd2653] <= 32'd1729;
		word[15'd2654] <= 32'd1730;
		word[15'd2655] <= 32'd1731;
		word[15'd2656] <= 32'd1732;
		word[15'd2657] <= 32'd1733;
		word[15'd2658] <= 32'd1734;
		word[15'd2659] <= 32'd1735;
		word[15'd2660] <= 32'd1736;
		word[15'd2661] <= 32'd1737;
		word[15'd2662] <= 32'd1738;
		word[15'd2663] <= 32'd1739;
		word[15'd2664] <= 32'd1740;
		word[15'd2665] <= 32'd1741;
		word[15'd2666] <= 32'd1742;
		word[15'd2667] <= 32'd1743;
		word[15'd2668] <= 32'd1744;
		word[15'd2669] <= 32'd1745;
		word[15'd2670] <= 32'd1746;
		word[15'd2671] <= 32'd1747;
		word[15'd2672] <= 32'd1748;
		word[15'd2673] <= 32'd1749;
		word[15'd2674] <= 32'd1750;
		word[15'd2675] <= 32'd1751;
		word[15'd2676] <= 32'd1752;
		word[15'd2677] <= 32'd1753;
		word[15'd2678] <= 32'd1754;
		word[15'd2679] <= 32'd1755;
		word[15'd2680] <= 32'd1756;
		word[15'd2681] <= 32'd1757;
		word[15'd2682] <= 32'd1758;
		word[15'd2683] <= 32'd1759;
		word[15'd2684] <= 32'd1760;
		word[15'd2685] <= 32'd1761;
		word[15'd2686] <= 32'd1762;
		word[15'd2687] <= 32'd1763;
		word[15'd2688] <= 32'd1764;
		word[15'd2689] <= 32'd1765;
		word[15'd2690] <= 32'd1766;
		word[15'd2691] <= 32'd1767;
		word[15'd2692] <= 32'd1768;
		word[15'd2693] <= 32'd1769;
		word[15'd2694] <= 32'd1770;
		word[15'd2695] <= 32'd1771;
		word[15'd2696] <= 32'd1772;
		word[15'd2697] <= 32'd1773;
		word[15'd2698] <= 32'd1774;
		word[15'd2699] <= 32'd1775;
		word[15'd2700] <= 32'd1776;
		word[15'd2701] <= 32'd1777;
		word[15'd2702] <= 32'd1778;
		word[15'd2703] <= 32'd1779;
		word[15'd2704] <= 32'd1780;
		word[15'd2705] <= 32'd1781;
		word[15'd2706] <= 32'd1782;
		word[15'd2707] <= 32'd1783;
		word[15'd2708] <= 32'd1784;
		word[15'd2709] <= 32'd1785;
		word[15'd2710] <= 32'd1786;
		word[15'd2711] <= 32'd1787;
		word[15'd2712] <= 32'd1788;
		word[15'd2713] <= 32'd1789;
		word[15'd2714] <= 32'd1790;
		word[15'd2715] <= 32'd1791;
		word[15'd2716] <= 32'd1792;
		word[15'd2717] <= 32'd1793;
		word[15'd2718] <= 32'd1794;
		word[15'd2719] <= 32'd1795;
		word[15'd2720] <= 32'd1796;
		word[15'd2721] <= 32'd1797;
		word[15'd2722] <= 32'd1798;
		word[15'd2723] <= 32'd1799;
		word[15'd2724] <= 32'd1800;
		word[15'd2725] <= 32'd1801;
		word[15'd2726] <= 32'd1802;
		word[15'd2727] <= 32'd1803;
		word[15'd2728] <= 32'd1804;
		word[15'd2729] <= 32'd1805;
		word[15'd2730] <= 32'd1806;
		word[15'd2731] <= 32'd1807;
		word[15'd2732] <= 32'd1808;
		word[15'd2733] <= 32'd1809;
		word[15'd2734] <= 32'd1810;
		word[15'd2735] <= 32'd1811;
		word[15'd2736] <= 32'd1812;
		word[15'd2737] <= 32'd1813;
		word[15'd2738] <= 32'd1814;
		word[15'd2739] <= 32'd1815;
		word[15'd2740] <= 32'd1816;
		word[15'd2741] <= 32'd1817;
		word[15'd2742] <= 32'd1818;
		word[15'd2743] <= 32'd1819;
		word[15'd2744] <= 32'd1820;
		word[15'd2745] <= 32'd1821;
		word[15'd2746] <= 32'd1822;
		word[15'd2747] <= 32'd1823;
		word[15'd2748] <= 32'd1824;
		word[15'd2749] <= 32'd1825;
		word[15'd2750] <= 32'd1826;
		word[15'd2751] <= 32'd1827;
		word[15'd2752] <= 32'd1828;
		word[15'd2753] <= 32'd1829;
		word[15'd2754] <= 32'd1830;
		word[15'd2755] <= 32'd1831;
		word[15'd2756] <= 32'd1832;
		word[15'd2757] <= 32'd1833;
		word[15'd2758] <= 32'd1834;
		word[15'd2759] <= 32'd1835;
		word[15'd2760] <= 32'd1836;
		word[15'd2761] <= 32'd1837;
		word[15'd2762] <= 32'd1838;
		word[15'd2763] <= 32'd1839;
		word[15'd2764] <= 32'd1840;
		word[15'd2765] <= 32'd1841;
		word[15'd2766] <= 32'd1842;
		word[15'd2767] <= 32'd1843;
		word[15'd2768] <= 32'd1844;
		word[15'd2769] <= 32'd1845;
		word[15'd2770] <= 32'd1846;
		word[15'd2771] <= 32'd1847;
		word[15'd2772] <= 32'd1848;
		word[15'd2773] <= 32'd1849;
		word[15'd2774] <= 32'd1850;
		word[15'd2775] <= 32'd1851;
		word[15'd2776] <= 32'd1852;
		word[15'd2777] <= 32'd1853;
		word[15'd2778] <= 32'd1854;
		word[15'd2779] <= 32'd1855;
		word[15'd2780] <= 32'd1856;
		word[15'd2781] <= 32'd1857;
		word[15'd2782] <= 32'd1858;
		word[15'd2783] <= 32'd1859;
		word[15'd2784] <= 32'd1860;
		word[15'd2785] <= 32'd1861;
		word[15'd2786] <= 32'd1862;
		word[15'd2787] <= 32'd1863;
		word[15'd2788] <= 32'd1864;
		word[15'd2789] <= 32'd1865;
		word[15'd2790] <= 32'd1866;
		word[15'd2791] <= 32'd1867;
		word[15'd2792] <= 32'd1868;
		word[15'd2793] <= 32'd1869;
		word[15'd2794] <= 32'd1870;
		word[15'd2795] <= 32'd1871;
		word[15'd2796] <= 32'd1872;
		word[15'd2797] <= 32'd1873;
		word[15'd2798] <= 32'd1874;
		word[15'd2799] <= 32'd1875;
		word[15'd2800] <= 32'd1876;
		word[15'd2801] <= 32'd1877;
		word[15'd2802] <= 32'd1878;
		word[15'd2803] <= 32'd1879;
		word[15'd2804] <= 32'd1880;
		word[15'd2805] <= 32'd1881;
		word[15'd2806] <= 32'd1882;
		word[15'd2807] <= 32'd1883;
		word[15'd2808] <= 32'd1884;
		word[15'd2809] <= 32'd1885;
		word[15'd2810] <= 32'd1886;
		word[15'd2811] <= 32'd1887;
		word[15'd2812] <= 32'd1888;
		word[15'd2813] <= 32'd1889;
		word[15'd2814] <= 32'd1890;
		word[15'd2815] <= 32'd1891;
		word[15'd2816] <= 32'd1892;
		word[15'd2817] <= 32'd1893;
		word[15'd2818] <= 32'd1894;
		word[15'd2819] <= 32'd1895;
		word[15'd2820] <= 32'd1896;
		word[15'd2821] <= 32'd1897;
		word[15'd2822] <= 32'd1898;
		word[15'd2823] <= 32'd1899;
		word[15'd2824] <= 32'd1900;
		word[15'd2825] <= 32'd1901;
		word[15'd2826] <= 32'd1902;
		word[15'd2827] <= 32'd1903;
		word[15'd2828] <= 32'd1904;
		word[15'd2829] <= 32'd1905;
		word[15'd2830] <= 32'd1906;
		word[15'd2831] <= 32'd1907;
		word[15'd2832] <= 32'd1908;
		word[15'd2833] <= 32'd1909;
		word[15'd2834] <= 32'd1910;
		word[15'd2835] <= 32'd1911;
		word[15'd2836] <= 32'd1912;
		word[15'd2837] <= 32'd1913;
		word[15'd2838] <= 32'd1914;
		word[15'd2839] <= 32'd1915;
		word[15'd2840] <= 32'd1916;
		word[15'd2841] <= 32'd1917;
		word[15'd2842] <= 32'd1918;
		word[15'd2843] <= 32'd1919;
		word[15'd2844] <= 32'd1920;
		word[15'd2845] <= 32'd1921;
		word[15'd2846] <= 32'd1922;
		word[15'd2847] <= 32'd1923;
		word[15'd2848] <= 32'd1924;
		word[15'd2849] <= 32'd1925;
		word[15'd2850] <= 32'd1926;
		word[15'd2851] <= 32'd1927;
		word[15'd2852] <= 32'd1928;
		word[15'd2853] <= 32'd1929;
		word[15'd2854] <= 32'd1930;
		word[15'd2855] <= 32'd1931;
		word[15'd2856] <= 32'd1932;
		word[15'd2857] <= 32'd1933;
		word[15'd2858] <= 32'd1934;
		word[15'd2859] <= 32'd1935;
		word[15'd2860] <= 32'd1936;
		word[15'd2861] <= 32'd1937;
		word[15'd2862] <= 32'd1938;
		word[15'd2863] <= 32'd1939;
		word[15'd2864] <= 32'd1940;
		word[15'd2865] <= 32'd1941;
		word[15'd2866] <= 32'd1942;
		word[15'd2867] <= 32'd1943;
		word[15'd2868] <= 32'd1944;
		word[15'd2869] <= 32'd1945;
		word[15'd2870] <= 32'd1946;
		word[15'd2871] <= 32'd1947;
		word[15'd2872] <= 32'd1948;
		word[15'd2873] <= 32'd1949;
		word[15'd2874] <= 32'd1950;
		word[15'd2875] <= 32'd1951;
		word[15'd2876] <= 32'd1952;
		word[15'd2877] <= 32'd1953;
		word[15'd2878] <= 32'd1954;
		word[15'd2879] <= 32'd1955;
		word[15'd2880] <= 32'd1956;
		word[15'd2881] <= 32'd1957;
		word[15'd2882] <= 32'd1958;
		word[15'd2883] <= 32'd1959;
		word[15'd2884] <= 32'd1960;
		word[15'd2885] <= 32'd1961;
		word[15'd2886] <= 32'd1962;
		word[15'd2887] <= 32'd1963;
		word[15'd2888] <= 32'd1964;
		word[15'd2889] <= 32'd1965;
		word[15'd2890] <= 32'd1966;
		word[15'd2891] <= 32'd1967;
		word[15'd2892] <= 32'd1968;
		word[15'd2893] <= 32'd1969;
		word[15'd2894] <= 32'd1970;
		word[15'd2895] <= 32'd1971;
		word[15'd2896] <= 32'd1972;
		word[15'd2897] <= 32'd1973;
		word[15'd2898] <= 32'd1974;
		word[15'd2899] <= 32'd1975;
		word[15'd2900] <= 32'd1976;
		word[15'd2901] <= 32'd1977;
		word[15'd2902] <= 32'd1978;
		word[15'd2903] <= 32'd1979;
		word[15'd2904] <= 32'd1980;
		word[15'd2905] <= 32'd1981;
		word[15'd2906] <= 32'd1982;
		word[15'd2907] <= 32'd1983;
		word[15'd2908] <= 32'd1984;
		word[15'd2909] <= 32'd1985;
		word[15'd2910] <= 32'd1986;
		word[15'd2911] <= 32'd1987;
		word[15'd2912] <= 32'd1988;
		word[15'd2913] <= 32'd1989;
		word[15'd2914] <= 32'd1990;
		word[15'd2915] <= 32'd1991;
		word[15'd2916] <= 32'd1992;
		word[15'd2917] <= 32'd1993;
		word[15'd2918] <= 32'd1994;
		word[15'd2919] <= 32'd1995;
		word[15'd2920] <= 32'd1996;
		word[15'd2921] <= 32'd1997;
		word[15'd2922] <= 32'd1998;
		word[15'd2923] <= 32'd1999;
		word[15'd2924] <= 32'd2000;
		word[15'd2925] <= 32'd2001;
		word[15'd2926] <= 32'd2002;
		word[15'd2927] <= 32'd2003;
		word[15'd2928] <= 32'd2004;
		word[15'd2929] <= 32'd2005;
		word[15'd2930] <= 32'd2006;
		word[15'd2931] <= 32'd2007;
		word[15'd2932] <= 32'd2008;
		word[15'd2933] <= 32'd2009;
		word[15'd2934] <= 32'd2010;
		word[15'd2935] <= 32'd2011;
		word[15'd2936] <= 32'd2012;
		word[15'd2937] <= 32'd2013;
		word[15'd2938] <= 32'd2014;
		word[15'd2939] <= 32'd2015;
		word[15'd2940] <= 32'd2016;
		word[15'd2941] <= 32'd2017;
		word[15'd2942] <= 32'd2018;
		word[15'd2943] <= 32'd2019;
		word[15'd2944] <= 32'd2020;
		word[15'd2945] <= 32'd2021;
		word[15'd2946] <= 32'd2022;
		word[15'd2947] <= 32'd2023;
		word[15'd2948] <= 32'd2024;
		word[15'd2949] <= 32'd2025;
		word[15'd2950] <= 32'd2026;
		word[15'd2951] <= 32'd2027;
		word[15'd2952] <= 32'd2028;
		word[15'd2953] <= 32'd2029;
		word[15'd2954] <= 32'd2030;
		word[15'd2955] <= 32'd2031;
		word[15'd2956] <= 32'd2032;
		word[15'd2957] <= 32'd2033;
		word[15'd2958] <= 32'd2034;
		word[15'd2959] <= 32'd2035;
		word[15'd2960] <= 32'd2036;
		word[15'd2961] <= 32'd2037;
		word[15'd2962] <= 32'd2038;
		word[15'd2963] <= 32'd2039;
		word[15'd2964] <= 32'd2040;
		word[15'd2965] <= 32'd2041;
		word[15'd2966] <= 32'd2042;
		word[15'd2967] <= 32'd2043;
		word[15'd2968] <= 32'd2044;
		word[15'd2969] <= 32'd2045;
		word[15'd2970] <= 32'd2046;
		word[15'd2971] <= 32'd2047;
		word[15'd2972] <= 32'd2048;
		word[15'd2973] <= 32'd2049;
		word[15'd2974] <= 32'd2050;
		word[15'd2975] <= 32'd2051;
		word[15'd2976] <= 32'd2052;
		word[15'd2977] <= 32'd2053;
		word[15'd2978] <= 32'd2054;
		word[15'd2979] <= 32'd2055;
		word[15'd2980] <= 32'd2056;
		word[15'd2981] <= 32'd2057;
		word[15'd2982] <= 32'd2058;
		word[15'd2983] <= 32'd2059;
		word[15'd2984] <= 32'd2060;
		word[15'd2985] <= 32'd2061;
		word[15'd2986] <= 32'd2062;
		word[15'd2987] <= 32'd2063;
		word[15'd2988] <= 32'd2064;
		word[15'd2989] <= 32'd2065;
		word[15'd2990] <= 32'd2066;
		word[15'd2991] <= 32'd2067;
		word[15'd2992] <= 32'd2068;
		word[15'd2993] <= 32'd2069;
		word[15'd2994] <= 32'd2070;
		word[15'd2995] <= 32'd2071;
		word[15'd2996] <= 32'd2072;
		word[15'd2997] <= 32'd2073;
		word[15'd2998] <= 32'd2074;
		word[15'd2999] <= 32'd2075;
		word[15'd3000] <= 32'd2076;
		word[15'd3001] <= 32'd2077;
		word[15'd3002] <= 32'd2078;
		word[15'd3003] <= 32'd2079;
		word[15'd3004] <= 32'd2080;
		word[15'd3005] <= 32'd2081;
		word[15'd3006] <= 32'd2082;
		word[15'd3007] <= 32'd2083;
		word[15'd3008] <= 32'd2084;
		word[15'd3009] <= 32'd2085;
		word[15'd3010] <= 32'd2086;
		word[15'd3011] <= 32'd2087;
		word[15'd3012] <= 32'd2088;
		word[15'd3013] <= 32'd2089;
		word[15'd3014] <= 32'd2090;
		word[15'd3015] <= 32'd2091;
		word[15'd3016] <= 32'd2092;
		word[15'd3017] <= 32'd2093;
		word[15'd3018] <= 32'd2094;
		word[15'd3019] <= 32'd2095;
		word[15'd3020] <= 32'd2096;
		word[15'd3021] <= 32'd2097;
		word[15'd3022] <= 32'd2098;
		word[15'd3023] <= 32'd2099;
		word[15'd3024] <= 32'd2100;
		word[15'd3025] <= 32'd2101;
		word[15'd3026] <= 32'd2102;
		word[15'd3027] <= 32'd2103;
		word[15'd3028] <= 32'd2104;
		word[15'd3029] <= 32'd2105;
		word[15'd3030] <= 32'd2106;
		word[15'd3031] <= 32'd2107;
		word[15'd3032] <= 32'd2108;
		word[15'd3033] <= 32'd2109;
		word[15'd3034] <= 32'd2110;
		word[15'd3035] <= 32'd2111;
		word[15'd3036] <= 32'd2112;
		word[15'd3037] <= 32'd2113;
		word[15'd3038] <= 32'd2114;
		word[15'd3039] <= 32'd2115;
		word[15'd3040] <= 32'd2116;
		word[15'd3041] <= 32'd2117;
		word[15'd3042] <= 32'd2118;
		word[15'd3043] <= 32'd2119;
		word[15'd3044] <= 32'd2120;
		word[15'd3045] <= 32'd2121;
		word[15'd3046] <= 32'd2122;
		word[15'd3047] <= 32'd2123;
		word[15'd3048] <= 32'd2124;
		word[15'd3049] <= 32'd2125;
		word[15'd3050] <= 32'd2126;
		word[15'd3051] <= 32'd2127;
		word[15'd3052] <= 32'd2128;
		word[15'd3053] <= 32'd2129;
		word[15'd3054] <= 32'd2130;
		word[15'd3055] <= 32'd2131;
		word[15'd3056] <= 32'd2132;
		word[15'd3057] <= 32'd2133;
		word[15'd3058] <= 32'd2134;
		word[15'd3059] <= 32'd2135;
		word[15'd3060] <= 32'd2136;
		word[15'd3061] <= 32'd2137;
		word[15'd3062] <= 32'd2138;
		word[15'd3063] <= 32'd2139;
		word[15'd3064] <= 32'd2140;
		word[15'd3065] <= 32'd2141;
		word[15'd3066] <= 32'd2142;
		word[15'd3067] <= 32'd2143;
		word[15'd3068] <= 32'd2144;
		word[15'd3069] <= 32'd2145;
		word[15'd3070] <= 32'd2146;
		word[15'd3071] <= 32'd2147;
		word[15'd3072] <= 32'd2148;
		word[15'd3073] <= 32'd2149;
		word[15'd3074] <= 32'd2150;
		word[15'd3075] <= 32'd2151;
		word[15'd3076] <= 32'd2152;
		word[15'd3077] <= 32'd2153;
		word[15'd3078] <= 32'd2154;
		word[15'd3079] <= 32'd2155;
		word[15'd3080] <= 32'd2156;
		word[15'd3081] <= 32'd2157;
		word[15'd3082] <= 32'd2158;
		word[15'd3083] <= 32'd2159;
		word[15'd3084] <= 32'd2160;
		word[15'd3085] <= 32'd2161;
		word[15'd3086] <= 32'd2162;
		word[15'd3087] <= 32'd2163;
		word[15'd3088] <= 32'd2164;
		word[15'd3089] <= 32'd2165;
		word[15'd3090] <= 32'd2166;
		word[15'd3091] <= 32'd2167;
		word[15'd3092] <= 32'd2168;
		word[15'd3093] <= 32'd2169;
		word[15'd3094] <= 32'd2170;
		word[15'd3095] <= 32'd2171;
		word[15'd3096] <= 32'd2172;
		word[15'd3097] <= 32'd2173;
		word[15'd3098] <= 32'd2174;
		word[15'd3099] <= 32'd2175;
		word[15'd3100] <= 32'd2176;
		word[15'd3101] <= 32'd2177;
		word[15'd3102] <= 32'd2178;
		word[15'd3103] <= 32'd2179;
		word[15'd3104] <= 32'd2180;
		word[15'd3105] <= 32'd2181;
		word[15'd3106] <= 32'd2182;
		word[15'd3107] <= 32'd2183;
		word[15'd3108] <= 32'd2184;
		word[15'd3109] <= 32'd2185;
		word[15'd3110] <= 32'd2186;
		word[15'd3111] <= 32'd2187;
		word[15'd3112] <= 32'd2188;
		word[15'd3113] <= 32'd2189;
		word[15'd3114] <= 32'd2190;
		word[15'd3115] <= 32'd2191;
		word[15'd3116] <= 32'd2192;
		word[15'd3117] <= 32'd2193;
		word[15'd3118] <= 32'd2194;
		word[15'd3119] <= 32'd2195;
		word[15'd3120] <= 32'd2196;
		word[15'd3121] <= 32'd2197;
		word[15'd3122] <= 32'd2198;
		word[15'd3123] <= 32'd2199;
		word[15'd3124] <= 32'd2200;
		word[15'd3125] <= 32'd2201;
		word[15'd3126] <= 32'd2202;
		word[15'd3127] <= 32'd2203;
		word[15'd3128] <= 32'd2204;
		word[15'd3129] <= 32'd2205;
		word[15'd3130] <= 32'd2206;
		word[15'd3131] <= 32'd2207;
		word[15'd3132] <= 32'd2208;
		word[15'd3133] <= 32'd2209;
		word[15'd3134] <= 32'd2210;
		word[15'd3135] <= 32'd2211;
		word[15'd3136] <= 32'd2212;
		word[15'd3137] <= 32'd2213;
		word[15'd3138] <= 32'd2214;
		word[15'd3139] <= 32'd2215;
		word[15'd3140] <= 32'd2216;
		word[15'd3141] <= 32'd2217;
		word[15'd3142] <= 32'd2218;
		word[15'd3143] <= 32'd2219;
		word[15'd3144] <= 32'd2220;
		word[15'd3145] <= 32'd2221;
		word[15'd3146] <= 32'd2222;
		word[15'd3147] <= 32'd2223;
		word[15'd3148] <= 32'd2224;
		word[15'd3149] <= 32'd2225;
		word[15'd3150] <= 32'd2226;
		word[15'd3151] <= 32'd2227;
		word[15'd3152] <= 32'd2228;
		word[15'd3153] <= 32'd2229;
		word[15'd3154] <= 32'd2230;
		word[15'd3155] <= 32'd2231;
		word[15'd3156] <= 32'd2232;
		word[15'd3157] <= 32'd2233;
		word[15'd3158] <= 32'd2234;
		word[15'd3159] <= 32'd2235;
		word[15'd3160] <= 32'd2236;
		word[15'd3161] <= 32'd2237;
		word[15'd3162] <= 32'd2238;
		word[15'd3163] <= 32'd2239;
		word[15'd3164] <= 32'd2240;
		word[15'd3165] <= 32'd2241;
		word[15'd3166] <= 32'd2242;
		word[15'd3167] <= 32'd2243;
		word[15'd3168] <= 32'd2244;
		word[15'd3169] <= 32'd2245;
		word[15'd3170] <= 32'd2246;
		word[15'd3171] <= 32'd2247;
		word[15'd3172] <= 32'd2248;
		word[15'd3173] <= 32'd2249;
		word[15'd3174] <= 32'd2250;
		word[15'd3175] <= 32'd2251;
		word[15'd3176] <= 32'd2252;
		word[15'd3177] <= 32'd2253;
		word[15'd3178] <= 32'd2254;
		word[15'd3179] <= 32'd2255;
		word[15'd3180] <= 32'd2256;
		word[15'd3181] <= 32'd2257;
		word[15'd3182] <= 32'd2258;
		word[15'd3183] <= 32'd2259;
		word[15'd3184] <= 32'd2260;
		word[15'd3185] <= 32'd2261;
		word[15'd3186] <= 32'd2262;
		word[15'd3187] <= 32'd2263;
		word[15'd3188] <= 32'd2264;
		word[15'd3189] <= 32'd2265;
		word[15'd3190] <= 32'd2266;
		word[15'd3191] <= 32'd2267;
		word[15'd3192] <= 32'd2268;
		word[15'd3193] <= 32'd2269;
		word[15'd3194] <= 32'd2270;
		word[15'd3195] <= 32'd2271;
		word[15'd3196] <= 32'd2272;
		word[15'd3197] <= 32'd2273;
		word[15'd3198] <= 32'd2274;
		word[15'd3199] <= 32'd2275;
		word[15'd3200] <= 32'd2276;
		word[15'd3201] <= 32'd2277;
		word[15'd3202] <= 32'd2278;
		word[15'd3203] <= 32'd2279;
		word[15'd3204] <= 32'd2280;
		word[15'd3205] <= 32'd2281;
		word[15'd3206] <= 32'd2282;
		word[15'd3207] <= 32'd2283;
		word[15'd3208] <= 32'd2284;
		word[15'd3209] <= 32'd2285;
		word[15'd3210] <= 32'd2286;
		word[15'd3211] <= 32'd2287;
		word[15'd3212] <= 32'd2288;
		word[15'd3213] <= 32'd2289;
		word[15'd3214] <= 32'd2290;
		word[15'd3215] <= 32'd2291;
		word[15'd3216] <= 32'd2292;
		word[15'd3217] <= 32'd2293;
		word[15'd3218] <= 32'd2294;
		word[15'd3219] <= 32'd2295;
		word[15'd3220] <= 32'd2296;
		word[15'd3221] <= 32'd2297;
		word[15'd3222] <= 32'd2298;
		word[15'd3223] <= 32'd2299;
		word[15'd3224] <= 32'd2300;
		word[15'd3225] <= 32'd2301;
		word[15'd3226] <= 32'd2302;
		word[15'd3227] <= 32'd2303;
		word[15'd3228] <= 32'd2304;
		word[15'd3229] <= 32'd2305;
		word[15'd3230] <= 32'd2306;
		word[15'd3231] <= 32'd2307;
		word[15'd3232] <= 32'd2308;
		word[15'd3233] <= 32'd2309;
		word[15'd3234] <= 32'd2310;
		word[15'd3235] <= 32'd2311;
		word[15'd3236] <= 32'd2312;
		word[15'd3237] <= 32'd2313;
		word[15'd3238] <= 32'd2314;
		word[15'd3239] <= 32'd2315;
		word[15'd3240] <= 32'd2316;
		word[15'd3241] <= 32'd2317;
		word[15'd3242] <= 32'd2318;
		word[15'd3243] <= 32'd2319;
		word[15'd3244] <= 32'd2320;
		word[15'd3245] <= 32'd2321;
		word[15'd3246] <= 32'd2322;
		word[15'd3247] <= 32'd2323;
		word[15'd3248] <= 32'd2324;
		word[15'd3249] <= 32'd2325;
		word[15'd3250] <= 32'd2326;
		word[15'd3251] <= 32'd2327;
		word[15'd3252] <= 32'd2328;
		word[15'd3253] <= 32'd2329;
		word[15'd3254] <= 32'd2330;
		word[15'd3255] <= 32'd2331;
		word[15'd3256] <= 32'd2332;
		word[15'd3257] <= 32'd2333;
		word[15'd3258] <= 32'd2334;
		word[15'd3259] <= 32'd2335;
		word[15'd3260] <= 32'd2336;
		word[15'd3261] <= 32'd2337;
		word[15'd3262] <= 32'd2338;
		word[15'd3263] <= 32'd2339;
		word[15'd3264] <= 32'd2340;
		word[15'd3265] <= 32'd2341;
		word[15'd3266] <= 32'd2342;
		word[15'd3267] <= 32'd2343;
		word[15'd3268] <= 32'd2344;
		word[15'd3269] <= 32'd2345;
		word[15'd3270] <= 32'd2346;
		word[15'd3271] <= 32'd2347;
		word[15'd3272] <= 32'd2348;
		word[15'd3273] <= 32'd2349;
		word[15'd3274] <= 32'd2350;
		word[15'd3275] <= 32'd2351;
		word[15'd3276] <= 32'd2352;
		word[15'd3277] <= 32'd2353;
		word[15'd3278] <= 32'd2354;
		word[15'd3279] <= 32'd2355;
		word[15'd3280] <= 32'd2356;
		word[15'd3281] <= 32'd2357;
		word[15'd3282] <= 32'd2358;
		word[15'd3283] <= 32'd2359;
		word[15'd3284] <= 32'd2360;
		word[15'd3285] <= 32'd2361;
		word[15'd3286] <= 32'd2362;
		word[15'd3287] <= 32'd2363;
		word[15'd3288] <= 32'd2364;
		word[15'd3289] <= 32'd2365;
		word[15'd3290] <= 32'd2366;
		word[15'd3291] <= 32'd2367;
		word[15'd3292] <= 32'd2368;
		word[15'd3293] <= 32'd2369;
		word[15'd3294] <= 32'd2370;
		word[15'd3295] <= 32'd2371;
		word[15'd3296] <= 32'd2372;
		word[15'd3297] <= 32'd2373;
		word[15'd3298] <= 32'd2374;
		word[15'd3299] <= 32'd2375;
		word[15'd3300] <= 32'd2376;
		word[15'd3301] <= 32'd2377;
		word[15'd3302] <= 32'd2378;
		word[15'd3303] <= 32'd2379;
		word[15'd3304] <= 32'd2380;
		word[15'd3305] <= 32'd2381;
		word[15'd3306] <= 32'd2382;
		word[15'd3307] <= 32'd2383;
		word[15'd3308] <= 32'd2384;
		word[15'd3309] <= 32'd2385;
		word[15'd3310] <= 32'd2386;
		word[15'd3311] <= 32'd2387;
		word[15'd3312] <= 32'd2388;
		word[15'd3313] <= 32'd2389;
		word[15'd3314] <= 32'd2390;
		word[15'd3315] <= 32'd2391;
		word[15'd3316] <= 32'd2392;
		word[15'd3317] <= 32'd2393;
		word[15'd3318] <= 32'd2394;
		word[15'd3319] <= 32'd2395;
		word[15'd3320] <= 32'd2396;
		word[15'd3321] <= 32'd2397;
		word[15'd3322] <= 32'd2398;
		word[15'd3323] <= 32'd2399;
		word[15'd3324] <= 32'd2400;
		word[15'd3325] <= 32'd2401;
		word[15'd3326] <= 32'd2402;
		word[15'd3327] <= 32'd2403;
		word[15'd3328] <= 32'd2404;
		word[15'd3329] <= 32'd2405;
		word[15'd3330] <= 32'd2406;
		word[15'd3331] <= 32'd2407;
		word[15'd3332] <= 32'd2408;
		word[15'd3333] <= 32'd2409;
		word[15'd3334] <= 32'd2410;
		word[15'd3335] <= 32'd2411;
		word[15'd3336] <= 32'd2412;
		word[15'd3337] <= 32'd2413;
		word[15'd3338] <= 32'd2414;
		word[15'd3339] <= 32'd2415;
		word[15'd3340] <= 32'd2416;
		word[15'd3341] <= 32'd2417;
		word[15'd3342] <= 32'd2418;
		word[15'd3343] <= 32'd2419;
		word[15'd3344] <= 32'd2420;
		word[15'd3345] <= 32'd2421;
		word[15'd3346] <= 32'd2422;
		word[15'd3347] <= 32'd2423;
		word[15'd3348] <= 32'd2424;
		word[15'd3349] <= 32'd2425;
		word[15'd3350] <= 32'd2426;
		word[15'd3351] <= 32'd2427;
		word[15'd3352] <= 32'd2428;
		word[15'd3353] <= 32'd2429;
		word[15'd3354] <= 32'd2430;
		word[15'd3355] <= 32'd2431;
		word[15'd3356] <= 32'd2432;
		word[15'd3357] <= 32'd2433;
		word[15'd3358] <= 32'd2434;
		word[15'd3359] <= 32'd2435;
		word[15'd3360] <= 32'd2436;
		word[15'd3361] <= 32'd2437;
		word[15'd3362] <= 32'd2438;
		word[15'd3363] <= 32'd2439;
		word[15'd3364] <= 32'd2440;
		word[15'd3365] <= 32'd2441;
		word[15'd3366] <= 32'd2442;
		word[15'd3367] <= 32'd2443;
		word[15'd3368] <= 32'd2444;
		word[15'd3369] <= 32'd2445;
		word[15'd3370] <= 32'd2446;
		word[15'd3371] <= 32'd2447;
		word[15'd3372] <= 32'd2448;
		word[15'd3373] <= 32'd2449;
		word[15'd3374] <= 32'd2450;
		word[15'd3375] <= 32'd2451;
		word[15'd3376] <= 32'd2452;
		word[15'd3377] <= 32'd2453;
		word[15'd3378] <= 32'd2454;
		word[15'd3379] <= 32'd2455;
		word[15'd3380] <= 32'd2456;
		word[15'd3381] <= 32'd2457;
		word[15'd3382] <= 32'd2458;
		word[15'd3383] <= 32'd2459;
		word[15'd3384] <= 32'd2460;
		word[15'd3385] <= 32'd2461;
		word[15'd3386] <= 32'd2462;
		word[15'd3387] <= 32'd2463;
		word[15'd3388] <= 32'd2464;
		word[15'd3389] <= 32'd2465;
		word[15'd3390] <= 32'd2466;
		word[15'd3391] <= 32'd2467;
		word[15'd3392] <= 32'd2468;
		word[15'd3393] <= 32'd2469;
		word[15'd3394] <= 32'd2470;
		word[15'd3395] <= 32'd2471;
		word[15'd3396] <= 32'd2472;
		word[15'd3397] <= 32'd2473;
		word[15'd3398] <= 32'd2474;
		word[15'd3399] <= 32'd2475;
		word[15'd3400] <= 32'd2476;
		word[15'd3401] <= 32'd2477;
		word[15'd3402] <= 32'd2478;
		word[15'd3403] <= 32'd2479;
		word[15'd3404] <= 32'd2480;
		word[15'd3405] <= 32'd2481;
		word[15'd3406] <= 32'd2482;
		word[15'd3407] <= 32'd2483;
		word[15'd3408] <= 32'd2484;
		word[15'd3409] <= 32'd2485;
		word[15'd3410] <= 32'd2486;
		word[15'd3411] <= 32'd2487;
		word[15'd3412] <= 32'd2488;
		word[15'd3413] <= 32'd2489;
		word[15'd3414] <= 32'd2490;
		word[15'd3415] <= 32'd2491;
		word[15'd3416] <= 32'd2492;
		word[15'd3417] <= 32'd2493;
		word[15'd3418] <= 32'd2494;
		word[15'd3419] <= 32'd2495;
		word[15'd3420] <= 32'd2496;
		word[15'd3421] <= 32'd2497;
		word[15'd3422] <= 32'd2498;
		word[15'd3423] <= 32'd2499;
		word[15'd3424] <= 32'd2500;
		word[15'd3425] <= 32'd2501;
		word[15'd3426] <= 32'd2502;
		word[15'd3427] <= 32'd2503;
		word[15'd3428] <= 32'd2504;
		word[15'd3429] <= 32'd2505;
		word[15'd3430] <= 32'd2506;
		word[15'd3431] <= 32'd2507;
		word[15'd3432] <= 32'd2508;
		word[15'd3433] <= 32'd2509;
		word[15'd3434] <= 32'd2510;
		word[15'd3435] <= 32'd2511;
		word[15'd3436] <= 32'd2512;
		word[15'd3437] <= 32'd2513;
		word[15'd3438] <= 32'd2514;
		word[15'd3439] <= 32'd2515;
		word[15'd3440] <= 32'd2516;
		word[15'd3441] <= 32'd2517;
		word[15'd3442] <= 32'd2518;
		word[15'd3443] <= 32'd2519;
		word[15'd3444] <= 32'd2520;
		word[15'd3445] <= 32'd2521;
		word[15'd3446] <= 32'd2522;
		word[15'd3447] <= 32'd2523;
		word[15'd3448] <= 32'd2524;
		word[15'd3449] <= 32'd2525;
		word[15'd3450] <= 32'd2526;
		word[15'd3451] <= 32'd2527;
		word[15'd3452] <= 32'd2528;
		word[15'd3453] <= 32'd2529;
		word[15'd3454] <= 32'd2530;
		word[15'd3455] <= 32'd2531;
		word[15'd3456] <= 32'd2532;
		word[15'd3457] <= 32'd2533;
		word[15'd3458] <= 32'd2534;
		word[15'd3459] <= 32'd2535;
		word[15'd3460] <= 32'd2536;
		word[15'd3461] <= 32'd2537;
		word[15'd3462] <= 32'd2538;
		word[15'd3463] <= 32'd2539;
		word[15'd3464] <= 32'd2540;
		word[15'd3465] <= 32'd2541;
		word[15'd3466] <= 32'd2542;
		word[15'd3467] <= 32'd2543;
		word[15'd3468] <= 32'd2544;
		word[15'd3469] <= 32'd2545;
		word[15'd3470] <= 32'd2546;
		word[15'd3471] <= 32'd2547;
		word[15'd3472] <= 32'd2548;
		word[15'd3473] <= 32'd2549;
		word[15'd3474] <= 32'd2550;
		word[15'd3475] <= 32'd2551;
		word[15'd3476] <= 32'd2552;
		word[15'd3477] <= 32'd2553;
		word[15'd3478] <= 32'd2554;
		word[15'd3479] <= 32'd2555;
		word[15'd3480] <= 32'd2556;
		word[15'd3481] <= 32'd2557;
		word[15'd3482] <= 32'd2558;
		word[15'd3483] <= 32'd2559;
		word[15'd3484] <= 32'd2560;
		word[15'd3485] <= 32'd2561;
		word[15'd3486] <= 32'd2562;
		word[15'd3487] <= 32'd2563;
		word[15'd3488] <= 32'd2564;
		word[15'd3489] <= 32'd2565;
		word[15'd3490] <= 32'd2566;
		word[15'd3491] <= 32'd2567;
		word[15'd3492] <= 32'd2568;
		word[15'd3493] <= 32'd2569;
		word[15'd3494] <= 32'd2570;
		word[15'd3495] <= 32'd2571;
		word[15'd3496] <= 32'd2572;
		word[15'd3497] <= 32'd2573;
		word[15'd3498] <= 32'd2574;
		word[15'd3499] <= 32'd2575;
		word[15'd3500] <= 32'd2576;
		word[15'd3501] <= 32'd2577;
		word[15'd3502] <= 32'd2578;
		word[15'd3503] <= 32'd2579;
		word[15'd3504] <= 32'd2580;
		word[15'd3505] <= 32'd2581;
		word[15'd3506] <= 32'd2582;
		word[15'd3507] <= 32'd2583;
		word[15'd3508] <= 32'd2584;
		word[15'd3509] <= 32'd2585;
		word[15'd3510] <= 32'd2586;
		word[15'd3511] <= 32'd2587;
		word[15'd3512] <= 32'd2588;
		word[15'd3513] <= 32'd2589;
		word[15'd3514] <= 32'd2590;
		word[15'd3515] <= 32'd2591;
		word[15'd3516] <= 32'd2592;
		word[15'd3517] <= 32'd2593;
		word[15'd3518] <= 32'd2594;
		word[15'd3519] <= 32'd2595;
		word[15'd3520] <= 32'd2596;
		word[15'd3521] <= 32'd2597;
		word[15'd3522] <= 32'd2598;
		word[15'd3523] <= 32'd2599;
		word[15'd3524] <= 32'd2600;
		word[15'd3525] <= 32'd2601;
		word[15'd3526] <= 32'd2602;
		word[15'd3527] <= 32'd2603;
		word[15'd3528] <= 32'd2604;
		word[15'd3529] <= 32'd2605;
		word[15'd3530] <= 32'd2606;
		word[15'd3531] <= 32'd2607;
		word[15'd3532] <= 32'd2608;
		word[15'd3533] <= 32'd2609;
		word[15'd3534] <= 32'd2610;
		word[15'd3535] <= 32'd2611;
		word[15'd3536] <= 32'd2612;
		word[15'd3537] <= 32'd2613;
		word[15'd3538] <= 32'd2614;
		word[15'd3539] <= 32'd2615;
		word[15'd3540] <= 32'd2616;
		word[15'd3541] <= 32'd2617;
		word[15'd3542] <= 32'd2618;
		word[15'd3543] <= 32'd2619;
		word[15'd3544] <= 32'd2620;
		word[15'd3545] <= 32'd2621;
		word[15'd3546] <= 32'd2622;
		word[15'd3547] <= 32'd2623;
		word[15'd3548] <= 32'd2624;
		word[15'd3549] <= 32'd2625;
		word[15'd3550] <= 32'd2626;
		word[15'd3551] <= 32'd2627;
		word[15'd3552] <= 32'd2628;
		word[15'd3553] <= 32'd2629;
		word[15'd3554] <= 32'd2630;
		word[15'd3555] <= 32'd2631;
		word[15'd3556] <= 32'd2632;
		word[15'd3557] <= 32'd2633;
		word[15'd3558] <= 32'd2634;
		word[15'd3559] <= 32'd2635;
		word[15'd3560] <= 32'd2636;
		word[15'd3561] <= 32'd2637;
		word[15'd3562] <= 32'd2638;
		word[15'd3563] <= 32'd2639;
		word[15'd3564] <= 32'd2640;
		word[15'd3565] <= 32'd2641;
		word[15'd3566] <= 32'd2642;
		word[15'd3567] <= 32'd2643;
		word[15'd3568] <= 32'd2644;
		word[15'd3569] <= 32'd2645;
		word[15'd3570] <= 32'd2646;
		word[15'd3571] <= 32'd2647;
		word[15'd3572] <= 32'd2648;
		word[15'd3573] <= 32'd2649;
		word[15'd3574] <= 32'd2650;
		word[15'd3575] <= 32'd2651;
		word[15'd3576] <= 32'd2652;
		word[15'd3577] <= 32'd2653;
		word[15'd3578] <= 32'd2654;
		word[15'd3579] <= 32'd2655;
		word[15'd3580] <= 32'd2656;
		word[15'd3581] <= 32'd2657;
		word[15'd3582] <= 32'd2658;
		word[15'd3583] <= 32'd2659;
		word[15'd3584] <= 32'd2660;
		word[15'd3585] <= 32'd2661;
		word[15'd3586] <= 32'd2662;
		word[15'd3587] <= 32'd2663;
		word[15'd3588] <= 32'd2664;
		word[15'd3589] <= 32'd2665;
		word[15'd3590] <= 32'd2666;
		word[15'd3591] <= 32'd2667;
		word[15'd3592] <= 32'd2668;
		word[15'd3593] <= 32'd2669;
		word[15'd3594] <= 32'd2670;
		word[15'd3595] <= 32'd2671;
		word[15'd3596] <= 32'd2672;
		word[15'd3597] <= 32'd2673;
		word[15'd3598] <= 32'd2674;
		word[15'd3599] <= 32'd2675;
		word[15'd3600] <= 32'd2676;
		word[15'd3601] <= 32'd2677;
		word[15'd3602] <= 32'd2678;
		word[15'd3603] <= 32'd2679;
		word[15'd3604] <= 32'd2680;
		word[15'd3605] <= 32'd2681;
		word[15'd3606] <= 32'd2682;
		word[15'd3607] <= 32'd2683;
		word[15'd3608] <= 32'd2684;
		word[15'd3609] <= 32'd2685;
		word[15'd3610] <= 32'd2686;
		word[15'd3611] <= 32'd2687;
		word[15'd3612] <= 32'd2688;
		word[15'd3613] <= 32'd2689;
		word[15'd3614] <= 32'd2690;
		word[15'd3615] <= 32'd2691;
		word[15'd3616] <= 32'd2692;
		word[15'd3617] <= 32'd2693;
		word[15'd3618] <= 32'd2694;
		word[15'd3619] <= 32'd2695;
		word[15'd3620] <= 32'd2696;
		word[15'd3621] <= 32'd2697;
		word[15'd3622] <= 32'd2698;
		word[15'd3623] <= 32'd2699;
		word[15'd3624] <= 32'd2700;
		word[15'd3625] <= 32'd2701;
		word[15'd3626] <= 32'd2702;
		word[15'd3627] <= 32'd2703;
		word[15'd3628] <= 32'd2704;
		word[15'd3629] <= 32'd2705;
		word[15'd3630] <= 32'd2706;
		word[15'd3631] <= 32'd2707;
		word[15'd3632] <= 32'd2708;
		word[15'd3633] <= 32'd2709;
		word[15'd3634] <= 32'd2710;
		word[15'd3635] <= 32'd2711;
		word[15'd3636] <= 32'd2712;
		word[15'd3637] <= 32'd2713;
		word[15'd3638] <= 32'd2714;
		word[15'd3639] <= 32'd2715;
		word[15'd3640] <= 32'd2716;
		word[15'd3641] <= 32'd2717;
		word[15'd3642] <= 32'd2718;
		word[15'd3643] <= 32'd2719;
		word[15'd3644] <= 32'd2720;
		word[15'd3645] <= 32'd2721;
		word[15'd3646] <= 32'd2722;
		word[15'd3647] <= 32'd2723;
		word[15'd3648] <= 32'd2724;
		word[15'd3649] <= 32'd2725;
		word[15'd3650] <= 32'd2726;
		word[15'd3651] <= 32'd2727;
		word[15'd3652] <= 32'd2728;
		word[15'd3653] <= 32'd2729;
		word[15'd3654] <= 32'd2730;
		word[15'd3655] <= 32'd2731;
		word[15'd3656] <= 32'd2732;
		word[15'd3657] <= 32'd2733;
		word[15'd3658] <= 32'd2734;
		word[15'd3659] <= 32'd2735;
		word[15'd3660] <= 32'd2736;
		word[15'd3661] <= 32'd2737;
		word[15'd3662] <= 32'd2738;
		word[15'd3663] <= 32'd2739;
		word[15'd3664] <= 32'd2740;
		word[15'd3665] <= 32'd2741;
		word[15'd3666] <= 32'd2742;
		word[15'd3667] <= 32'd2743;
		word[15'd3668] <= 32'd2744;
		word[15'd3669] <= 32'd2745;
		word[15'd3670] <= 32'd2746;
		word[15'd3671] <= 32'd2747;
		word[15'd3672] <= 32'd2748;
		word[15'd3673] <= 32'd2749;
		word[15'd3674] <= 32'd2750;
		word[15'd3675] <= 32'd2751;
		word[15'd3676] <= 32'd2752;
		word[15'd3677] <= 32'd2753;
		word[15'd3678] <= 32'd2754;
		word[15'd3679] <= 32'd2755;
		word[15'd3680] <= 32'd2756;
		word[15'd3681] <= 32'd2757;
		word[15'd3682] <= 32'd2758;
		word[15'd3683] <= 32'd2759;
		word[15'd3684] <= 32'd2760;
		word[15'd3685] <= 32'd2761;
		word[15'd3686] <= 32'd2762;
		word[15'd3687] <= 32'd2763;
		word[15'd3688] <= 32'd2764;
		word[15'd3689] <= 32'd2765;
		word[15'd3690] <= 32'd2766;
		word[15'd3691] <= 32'd2767;
		word[15'd3692] <= 32'd2768;
		word[15'd3693] <= 32'd2769;
		word[15'd3694] <= 32'd2770;
		word[15'd3695] <= 32'd2771;
		word[15'd3696] <= 32'd2772;
		word[15'd3697] <= 32'd2773;
		word[15'd3698] <= 32'd2774;
		word[15'd3699] <= 32'd2775;
		word[15'd3700] <= 32'd2776;
		word[15'd3701] <= 32'd2777;
		word[15'd3702] <= 32'd2778;
		word[15'd3703] <= 32'd2779;
		word[15'd3704] <= 32'd2780;
		word[15'd3705] <= 32'd2781;
		word[15'd3706] <= 32'd2782;
		word[15'd3707] <= 32'd2783;
		word[15'd3708] <= 32'd2784;
		word[15'd3709] <= 32'd2785;
		word[15'd3710] <= 32'd2786;
		word[15'd3711] <= 32'd2787;
		word[15'd3712] <= 32'd2788;
		word[15'd3713] <= 32'd2789;
		word[15'd3714] <= 32'd2790;
		word[15'd3715] <= 32'd2791;
		word[15'd3716] <= 32'd2792;
		word[15'd3717] <= 32'd2793;
		word[15'd3718] <= 32'd2794;
		word[15'd3719] <= 32'd2795;
		word[15'd3720] <= 32'd2796;
		word[15'd3721] <= 32'd2797;
		word[15'd3722] <= 32'd2798;
		word[15'd3723] <= 32'd2799;
		word[15'd3724] <= 32'd2800;
		word[15'd3725] <= 32'd2801;
		word[15'd3726] <= 32'd2802;
		word[15'd3727] <= 32'd2803;
		word[15'd3728] <= 32'd2804;
		word[15'd3729] <= 32'd2805;
		word[15'd3730] <= 32'd2806;
		word[15'd3731] <= 32'd2807;
		word[15'd3732] <= 32'd2808;
		word[15'd3733] <= 32'd2809;
		word[15'd3734] <= 32'd2810;
		word[15'd3735] <= 32'd2811;
		word[15'd3736] <= 32'd2812;
		word[15'd3737] <= 32'd2813;
		word[15'd3738] <= 32'd2814;
		word[15'd3739] <= 32'd2815;
		word[15'd3740] <= 32'd2816;
		word[15'd3741] <= 32'd2817;
		word[15'd3742] <= 32'd2818;
		word[15'd3743] <= 32'd2819;
		word[15'd3744] <= 32'd2820;
		word[15'd3745] <= 32'd2821;
		word[15'd3746] <= 32'd2822;
		word[15'd3747] <= 32'd2823;
		word[15'd3748] <= 32'd2824;
		word[15'd3749] <= 32'd2825;
		word[15'd3750] <= 32'd2826;
		word[15'd3751] <= 32'd2827;
		word[15'd3752] <= 32'd2828;
		word[15'd3753] <= 32'd2829;
		word[15'd3754] <= 32'd2830;
		word[15'd3755] <= 32'd2831;
		word[15'd3756] <= 32'd2832;
		word[15'd3757] <= 32'd2833;
		word[15'd3758] <= 32'd2834;
		word[15'd3759] <= 32'd2835;
		word[15'd3760] <= 32'd2836;
		word[15'd3761] <= 32'd2837;
		word[15'd3762] <= 32'd2838;
		word[15'd3763] <= 32'd2839;
		word[15'd3764] <= 32'd2840;
		word[15'd3765] <= 32'd2841;
		word[15'd3766] <= 32'd2842;
		word[15'd3767] <= 32'd2843;
		word[15'd3768] <= 32'd2844;
		word[15'd3769] <= 32'd2845;
		word[15'd3770] <= 32'd2846;
		word[15'd3771] <= 32'd2847;
		word[15'd3772] <= 32'd2848;
		word[15'd3773] <= 32'd2849;
		word[15'd3774] <= 32'd2850;
		word[15'd3775] <= 32'd2851;
		word[15'd3776] <= 32'd2852;
		word[15'd3777] <= 32'd2853;
		word[15'd3778] <= 32'd2854;
		word[15'd3779] <= 32'd2855;
		word[15'd3780] <= 32'd2856;
		word[15'd3781] <= 32'd2857;
		word[15'd3782] <= 32'd2858;
		word[15'd3783] <= 32'd2859;
		word[15'd3784] <= 32'd2860;
		word[15'd3785] <= 32'd2861;
		word[15'd3786] <= 32'd2862;
		word[15'd3787] <= 32'd2863;
		word[15'd3788] <= 32'd2864;
		word[15'd3789] <= 32'd2865;
		word[15'd3790] <= 32'd2866;
		word[15'd3791] <= 32'd2867;
		word[15'd3792] <= 32'd2868;
		word[15'd3793] <= 32'd2869;
		word[15'd3794] <= 32'd2870;
		word[15'd3795] <= 32'd2871;
		word[15'd3796] <= 32'd2872;
		word[15'd3797] <= 32'd2873;
		word[15'd3798] <= 32'd2874;
		word[15'd3799] <= 32'd2875;
		word[15'd3800] <= 32'd2876;
		word[15'd3801] <= 32'd2877;
		word[15'd3802] <= 32'd2878;
		word[15'd3803] <= 32'd2879;
		word[15'd3804] <= 32'd2880;
		word[15'd3805] <= 32'd2881;
		word[15'd3806] <= 32'd2882;
		word[15'd3807] <= 32'd2883;
		word[15'd3808] <= 32'd2884;
		word[15'd3809] <= 32'd2885;
		word[15'd3810] <= 32'd2886;
		word[15'd3811] <= 32'd2887;
		word[15'd3812] <= 32'd2888;
		word[15'd3813] <= 32'd2889;
		word[15'd3814] <= 32'd2890;
		word[15'd3815] <= 32'd2891;
		word[15'd3816] <= 32'd2892;
		word[15'd3817] <= 32'd2893;
		word[15'd3818] <= 32'd2894;
		word[15'd3819] <= 32'd2895;
		word[15'd3820] <= 32'd2896;
		word[15'd3821] <= 32'd2897;
		word[15'd3822] <= 32'd2898;
		word[15'd3823] <= 32'd2899;
		word[15'd3824] <= 32'd2900;
		word[15'd3825] <= 32'd2901;
		word[15'd3826] <= 32'd2902;
		word[15'd3827] <= 32'd2903;
		word[15'd3828] <= 32'd2904;
		word[15'd3829] <= 32'd2905;
		word[15'd3830] <= 32'd2906;
		word[15'd3831] <= 32'd2907;
		word[15'd3832] <= 32'd2908;
		word[15'd3833] <= 32'd2909;
		word[15'd3834] <= 32'd2910;
		word[15'd3835] <= 32'd2911;
		word[15'd3836] <= 32'd2912;
		word[15'd3837] <= 32'd2913;
		word[15'd3838] <= 32'd2914;
		word[15'd3839] <= 32'd2915;
		word[15'd3840] <= 32'd2916;
		word[15'd3841] <= 32'd2917;
		word[15'd3842] <= 32'd2918;
		word[15'd3843] <= 32'd2919;
		word[15'd3844] <= 32'd2920;
		word[15'd3845] <= 32'd2921;
		word[15'd3846] <= 32'd2922;
		word[15'd3847] <= 32'd2923;
		word[15'd3848] <= 32'd2924;
		word[15'd3849] <= 32'd2925;
		word[15'd3850] <= 32'd2926;
		word[15'd3851] <= 32'd2927;
		word[15'd3852] <= 32'd2928;
		word[15'd3853] <= 32'd2929;
		word[15'd3854] <= 32'd2930;
		word[15'd3855] <= 32'd2931;
		word[15'd3856] <= 32'd2932;
		word[15'd3857] <= 32'd2933;
		word[15'd3858] <= 32'd2934;
		word[15'd3859] <= 32'd2935;
		word[15'd3860] <= 32'd2936;
		word[15'd3861] <= 32'd2937;
		word[15'd3862] <= 32'd2938;
		word[15'd3863] <= 32'd2939;
		word[15'd3864] <= 32'd2940;
		word[15'd3865] <= 32'd2941;
		word[15'd3866] <= 32'd2942;
		word[15'd3867] <= 32'd2943;
		word[15'd3868] <= 32'd2944;
		word[15'd3869] <= 32'd2945;
		word[15'd3870] <= 32'd2946;
		word[15'd3871] <= 32'd2947;
		word[15'd3872] <= 32'd2948;
		word[15'd3873] <= 32'd2949;
		word[15'd3874] <= 32'd2950;
		word[15'd3875] <= 32'd2951;
		word[15'd3876] <= 32'd2952;
		word[15'd3877] <= 32'd2953;
		word[15'd3878] <= 32'd2954;
		word[15'd3879] <= 32'd2955;
		word[15'd3880] <= 32'd2956;
		word[15'd3881] <= 32'd2957;
		word[15'd3882] <= 32'd2958;
		word[15'd3883] <= 32'd2959;
		word[15'd3884] <= 32'd2960;
		word[15'd3885] <= 32'd2961;
		word[15'd3886] <= 32'd2962;
		word[15'd3887] <= 32'd2963;
		word[15'd3888] <= 32'd2964;
		word[15'd3889] <= 32'd2965;
		word[15'd3890] <= 32'd2966;
		word[15'd3891] <= 32'd2967;
		word[15'd3892] <= 32'd2968;
		word[15'd3893] <= 32'd2969;
		word[15'd3894] <= 32'd2970;
		word[15'd3895] <= 32'd2971;
		word[15'd3896] <= 32'd2972;
		word[15'd3897] <= 32'd2973;
		word[15'd3898] <= 32'd2974;
		word[15'd3899] <= 32'd2975;
		word[15'd3900] <= 32'd2976;
		word[15'd3901] <= 32'd2977;
		word[15'd3902] <= 32'd2978;
		word[15'd3903] <= 32'd2979;
		word[15'd3904] <= 32'd2980;
		word[15'd3905] <= 32'd2981;
		word[15'd3906] <= 32'd2982;
		word[15'd3907] <= 32'd2983;
		word[15'd3908] <= 32'd2984;
		word[15'd3909] <= 32'd2985;
		word[15'd3910] <= 32'd2986;
		word[15'd3911] <= 32'd2987;
		word[15'd3912] <= 32'd2988;
		word[15'd3913] <= 32'd2989;
		word[15'd3914] <= 32'd2990;
		word[15'd3915] <= 32'd2991;
		word[15'd3916] <= 32'd2992;
		word[15'd3917] <= 32'd2993;
		word[15'd3918] <= 32'd2994;
		word[15'd3919] <= 32'd2995;
		word[15'd3920] <= 32'd2996;
		word[15'd3921] <= 32'd2997;
		word[15'd3922] <= 32'd2998;
		word[15'd3923] <= 32'd2999;
		word[15'd3924] <= 32'd3000;
		word[15'd3925] <= 32'd3001;
		word[15'd3926] <= 32'd3002;
		word[15'd3927] <= 32'd3003;
		word[15'd3928] <= 32'd3004;
		word[15'd3929] <= 32'd3005;
		word[15'd3930] <= 32'd3006;
		word[15'd3931] <= 32'd3007;
		word[15'd3932] <= 32'd3008;
		word[15'd3933] <= 32'd3009;
		word[15'd3934] <= 32'd3010;
		word[15'd3935] <= 32'd3011;
		word[15'd3936] <= 32'd3012;
		word[15'd3937] <= 32'd3013;
		word[15'd3938] <= 32'd3014;
		word[15'd3939] <= 32'd3015;
		word[15'd3940] <= 32'd3016;
		word[15'd3941] <= 32'd3017;
		word[15'd3942] <= 32'd3018;
		word[15'd3943] <= 32'd3019;
		word[15'd3944] <= 32'd3020;
		word[15'd3945] <= 32'd3021;
		word[15'd3946] <= 32'd3022;
		word[15'd3947] <= 32'd3023;
		word[15'd3948] <= 32'd3024;
		word[15'd3949] <= 32'd3025;
		word[15'd3950] <= 32'd3026;
		word[15'd3951] <= 32'd3027;
		word[15'd3952] <= 32'd3028;
		word[15'd3953] <= 32'd3029;
		word[15'd3954] <= 32'd3030;
		word[15'd3955] <= 32'd3031;
		word[15'd3956] <= 32'd3032;
		word[15'd3957] <= 32'd3033;
		word[15'd3958] <= 32'd3034;
		word[15'd3959] <= 32'd3035;
		word[15'd3960] <= 32'd3036;
		word[15'd3961] <= 32'd3037;
		word[15'd3962] <= 32'd3038;
		word[15'd3963] <= 32'd3039;
		word[15'd3964] <= 32'd3040;
		word[15'd3965] <= 32'd3041;
		word[15'd3966] <= 32'd3042;
		word[15'd3967] <= 32'd3043;
		word[15'd3968] <= 32'd3044;
		word[15'd3969] <= 32'd3045;
		word[15'd3970] <= 32'd3046;
		word[15'd3971] <= 32'd3047;
		word[15'd3972] <= 32'd3048;
		word[15'd3973] <= 32'd3049;
		word[15'd3974] <= 32'd3050;
		word[15'd3975] <= 32'd3051;
		word[15'd3976] <= 32'd3052;
		word[15'd3977] <= 32'd3053;
		word[15'd3978] <= 32'd3054;
		word[15'd3979] <= 32'd3055;
		word[15'd3980] <= 32'd3056;
		word[15'd3981] <= 32'd3057;
		word[15'd3982] <= 32'd3058;
		word[15'd3983] <= 32'd3059;
		word[15'd3984] <= 32'd3060;
		word[15'd3985] <= 32'd3061;
		word[15'd3986] <= 32'd3062;
		word[15'd3987] <= 32'd3063;
		word[15'd3988] <= 32'd3064;
		word[15'd3989] <= 32'd3065;
		word[15'd3990] <= 32'd3066;
		word[15'd3991] <= 32'd3067;
		word[15'd3992] <= 32'd3068;
		word[15'd3993] <= 32'd3069;
		word[15'd3994] <= 32'd3070;
		word[15'd3995] <= 32'd3071;
		word[15'd3996] <= 32'd3072;
		word[15'd3997] <= 32'd3073;
		word[15'd3998] <= 32'd3074;
		word[15'd3999] <= 32'd3075;
		word[15'd4000] <= 32'd3076;
		word[15'd4001] <= 32'd3077;
		word[15'd4002] <= 32'd3078;
		word[15'd4003] <= 32'd3079;
		word[15'd4004] <= 32'd3080;
		word[15'd4005] <= 32'd3081;
		word[15'd4006] <= 32'd3082;
		word[15'd4007] <= 32'd3083;
		word[15'd4008] <= 32'd3084;
		word[15'd4009] <= 32'd3085;
		word[15'd4010] <= 32'd3086;
		word[15'd4011] <= 32'd3087;
		word[15'd4012] <= 32'd3088;
		word[15'd4013] <= 32'd3089;
		word[15'd4014] <= 32'd3090;
		word[15'd4015] <= 32'd3091;
		word[15'd4016] <= 32'd3092;
		word[15'd4017] <= 32'd3093;
		word[15'd4018] <= 32'd3094;
		word[15'd4019] <= 32'd3095;
		word[15'd4020] <= 32'd3096;
		word[15'd4021] <= 32'd3097;
		word[15'd4022] <= 32'd3098;
		word[15'd4023] <= 32'd3099;
		word[15'd4024] <= 32'd3100;
		word[15'd4025] <= 32'd3101;
		word[15'd4026] <= 32'd3102;
		word[15'd4027] <= 32'd3103;
		word[15'd4028] <= 32'd3104;
		word[15'd4029] <= 32'd3105;
		word[15'd4030] <= 32'd3106;
		word[15'd4031] <= 32'd3107;
		word[15'd4032] <= 32'd3108;
		word[15'd4033] <= 32'd3109;
		word[15'd4034] <= 32'd3110;
		word[15'd4035] <= 32'd3111;
		word[15'd4036] <= 32'd3112;
		word[15'd4037] <= 32'd3113;
		word[15'd4038] <= 32'd3114;
		word[15'd4039] <= 32'd3115;
		word[15'd4040] <= 32'd3116;
		word[15'd4041] <= 32'd3117;
		word[15'd4042] <= 32'd3118;
		word[15'd4043] <= 32'd3119;
		word[15'd4044] <= 32'd3120;
		word[15'd4045] <= 32'd3121;
		word[15'd4046] <= 32'd3122;
		word[15'd4047] <= 32'd3123;
		word[15'd4048] <= 32'd3124;
		word[15'd4049] <= 32'd3125;
		word[15'd4050] <= 32'd3126;
		word[15'd4051] <= 32'd3127;
		word[15'd4052] <= 32'd3128;
		word[15'd4053] <= 32'd3129;
		word[15'd4054] <= 32'd3130;
		word[15'd4055] <= 32'd3131;
		word[15'd4056] <= 32'd3132;
		word[15'd4057] <= 32'd3133;
		word[15'd4058] <= 32'd3134;
		word[15'd4059] <= 32'd3135;
		word[15'd4060] <= 32'd3136;
		word[15'd4061] <= 32'd3137;
		word[15'd4062] <= 32'd3138;
		word[15'd4063] <= 32'd3139;
		word[15'd4064] <= 32'd3140;
		word[15'd4065] <= 32'd3141;
		word[15'd4066] <= 32'd3142;
		word[15'd4067] <= 32'd3143;
		word[15'd4068] <= 32'd3144;
		word[15'd4069] <= 32'd3145;
		word[15'd4070] <= 32'd3146;
		word[15'd4071] <= 32'd3147;
		word[15'd4072] <= 32'd3148;
		word[15'd4073] <= 32'd3149;
		word[15'd4074] <= 32'd3150;
		word[15'd4075] <= 32'd3151;
		word[15'd4076] <= 32'd3152;
		word[15'd4077] <= 32'd3153;
		word[15'd4078] <= 32'd3154;
		word[15'd4079] <= 32'd3155;
		word[15'd4080] <= 32'd3156;
		word[15'd4081] <= 32'd3157;
		word[15'd4082] <= 32'd3158;
		word[15'd4083] <= 32'd3159;
		word[15'd4084] <= 32'd3160;
		word[15'd4085] <= 32'd3161;
		word[15'd4086] <= 32'd3162;
		word[15'd4087] <= 32'd3163;
		word[15'd4088] <= 32'd3164;
		word[15'd4089] <= 32'd3165;
		word[15'd4090] <= 32'd3166;
		word[15'd4091] <= 32'd3167;
		word[15'd4092] <= 32'd3168;
		word[15'd4093] <= 32'd3169;
		word[15'd4094] <= 32'd3170;
		word[15'd4095] <= 32'd3171;
		word[15'd4096] <= 32'd3172;
		word[15'd4097] <= 32'd3173;
		word[15'd4098] <= 32'd3174;
		word[15'd4099] <= 32'd3175;
		word[15'd4100] <= 32'd3176;
		word[15'd4101] <= 32'd3177;
		word[15'd4102] <= 32'd3178;
		word[15'd4103] <= 32'd3179;
		word[15'd4104] <= 32'd3180;
		word[15'd4105] <= 32'd3181;
		word[15'd4106] <= 32'd3182;
		word[15'd4107] <= 32'd3183;
		word[15'd4108] <= 32'd3184;
		word[15'd4109] <= 32'd3185;
		word[15'd4110] <= 32'd3186;
		word[15'd4111] <= 32'd3187;
		word[15'd4112] <= 32'd3188;
		word[15'd4113] <= 32'd3189;
		word[15'd4114] <= 32'd3190;
		word[15'd4115] <= 32'd3191;
		word[15'd4116] <= 32'd3192;
		word[15'd4117] <= 32'd3193;
		word[15'd4118] <= 32'd3194;
		word[15'd4119] <= 32'd3195;
		word[15'd4120] <= 32'd3196;
		word[15'd4121] <= 32'd3197;
		word[15'd4122] <= 32'd3198;
		word[15'd4123] <= 32'd3199;
		word[15'd4124] <= 32'd3200;
		word[15'd4125] <= 32'd3201;
		word[15'd4126] <= 32'd3202;
		word[15'd4127] <= 32'd3203;
		word[15'd4128] <= 32'd3204;
		word[15'd4129] <= 32'd3205;
		word[15'd4130] <= 32'd3206;
		word[15'd4131] <= 32'd3207;
		word[15'd4132] <= 32'd3208;
		word[15'd4133] <= 32'd3209;
		word[15'd4134] <= 32'd3210;
		word[15'd4135] <= 32'd3211;
		word[15'd4136] <= 32'd3212;
		word[15'd4137] <= 32'd3213;
		word[15'd4138] <= 32'd3214;
		word[15'd4139] <= 32'd3215;
		word[15'd4140] <= 32'd3216;
		word[15'd4141] <= 32'd3217;
		word[15'd4142] <= 32'd3218;
		word[15'd4143] <= 32'd3219;
		word[15'd4144] <= 32'd3220;
		word[15'd4145] <= 32'd3221;
		word[15'd4146] <= 32'd3222;
		word[15'd4147] <= 32'd3223;
		word[15'd4148] <= 32'd3224;
		word[15'd4149] <= 32'd3225;
		word[15'd4150] <= 32'd3226;
		word[15'd4151] <= 32'd3227;
		word[15'd4152] <= 32'd3228;
		word[15'd4153] <= 32'd3229;
		word[15'd4154] <= 32'd3230;
		word[15'd4155] <= 32'd3231;
		word[15'd4156] <= 32'd3232;
		word[15'd4157] <= 32'd3233;
		word[15'd4158] <= 32'd3234;
		word[15'd4159] <= 32'd3235;
		word[15'd4160] <= 32'd3236;
		word[15'd4161] <= 32'd3237;
		word[15'd4162] <= 32'd3238;
		word[15'd4163] <= 32'd3239;
		word[15'd4164] <= 32'd3240;
		word[15'd4165] <= 32'd3241;
		word[15'd4166] <= 32'd3242;
		word[15'd4167] <= 32'd3243;
		word[15'd4168] <= 32'd3244;
		word[15'd4169] <= 32'd3245;
		word[15'd4170] <= 32'd3246;
		word[15'd4171] <= 32'd3247;
		word[15'd4172] <= 32'd3248;
		word[15'd4173] <= 32'd3249;
		word[15'd4174] <= 32'd3250;
		word[15'd4175] <= 32'd3251;
		word[15'd4176] <= 32'd3252;
		word[15'd4177] <= 32'd3253;
		word[15'd4178] <= 32'd3254;
		word[15'd4179] <= 32'd3255;
		word[15'd4180] <= 32'd3256;
		word[15'd4181] <= 32'd3257;
		word[15'd4182] <= 32'd3258;
		word[15'd4183] <= 32'd3259;
		word[15'd4184] <= 32'd3260;
		word[15'd4185] <= 32'd3261;
		word[15'd4186] <= 32'd3262;
		word[15'd4187] <= 32'd3263;
		word[15'd4188] <= 32'd3264;
		word[15'd4189] <= 32'd3265;
		word[15'd4190] <= 32'd3266;
		word[15'd4191] <= 32'd3267;
		word[15'd4192] <= 32'd3268;
		word[15'd4193] <= 32'd3269;
		word[15'd4194] <= 32'd3270;
		word[15'd4195] <= 32'd3271;
		word[15'd4196] <= 32'd3272;
		word[15'd4197] <= 32'd3273;
		word[15'd4198] <= 32'd3274;
		word[15'd4199] <= 32'd3275;
		word[15'd4200] <= 32'd3276;
		word[15'd4201] <= 32'd3277;
		word[15'd4202] <= 32'd3278;
		word[15'd4203] <= 32'd3279;
		word[15'd4204] <= 32'd3280;
		word[15'd4205] <= 32'd3281;
		word[15'd4206] <= 32'd3282;
		word[15'd4207] <= 32'd3283;
		word[15'd4208] <= 32'd3284;
		word[15'd4209] <= 32'd3285;
		word[15'd4210] <= 32'd3286;
		word[15'd4211] <= 32'd3287;
		word[15'd4212] <= 32'd3288;
		word[15'd4213] <= 32'd3289;
		word[15'd4214] <= 32'd3290;
		word[15'd4215] <= 32'd3291;
		word[15'd4216] <= 32'd3292;
		word[15'd4217] <= 32'd3293;
		word[15'd4218] <= 32'd3294;
		word[15'd4219] <= 32'd3295;
		word[15'd4220] <= 32'd3296;
		word[15'd4221] <= 32'd3297;
		word[15'd4222] <= 32'd3298;
		word[15'd4223] <= 32'd3299;
		word[15'd4224] <= 32'd3300;
		word[15'd4225] <= 32'd3301;
		word[15'd4226] <= 32'd3302;
		word[15'd4227] <= 32'd3303;
		word[15'd4228] <= 32'd3304;
		word[15'd4229] <= 32'd3305;
		word[15'd4230] <= 32'd3306;
		word[15'd4231] <= 32'd3307;
		word[15'd4232] <= 32'd3308;
		word[15'd4233] <= 32'd3309;
		word[15'd4234] <= 32'd3310;
		word[15'd4235] <= 32'd3311;
		word[15'd4236] <= 32'd3312;
		word[15'd4237] <= 32'd3313;
		word[15'd4238] <= 32'd3314;
		word[15'd4239] <= 32'd3315;
		word[15'd4240] <= 32'd3316;
		word[15'd4241] <= 32'd3317;
		word[15'd4242] <= 32'd3318;
		word[15'd4243] <= 32'd3319;
		word[15'd4244] <= 32'd3320;
		word[15'd4245] <= 32'd3321;
		word[15'd4246] <= 32'd3322;
		word[15'd4247] <= 32'd3323;
		word[15'd4248] <= 32'd3324;
		word[15'd4249] <= 32'd3325;
		word[15'd4250] <= 32'd3326;
		word[15'd4251] <= 32'd3327;
		word[15'd4252] <= 32'd3328;
		word[15'd4253] <= 32'd3329;
		word[15'd4254] <= 32'd3330;
		word[15'd4255] <= 32'd3331;
		word[15'd4256] <= 32'd3332;
		word[15'd4257] <= 32'd3333;
		word[15'd4258] <= 32'd3334;
		word[15'd4259] <= 32'd3335;
		word[15'd4260] <= 32'd3336;
		word[15'd4261] <= 32'd3337;
		word[15'd4262] <= 32'd3338;
		word[15'd4263] <= 32'd3339;
		word[15'd4264] <= 32'd3340;
		word[15'd4265] <= 32'd3341;
		word[15'd4266] <= 32'd3342;
		word[15'd4267] <= 32'd3343;
		word[15'd4268] <= 32'd3344;
		word[15'd4269] <= 32'd3345;
		word[15'd4270] <= 32'd3346;
		word[15'd4271] <= 32'd3347;
		word[15'd4272] <= 32'd3348;
		word[15'd4273] <= 32'd3349;
		word[15'd4274] <= 32'd3350;
		word[15'd4275] <= 32'd3351;
		word[15'd4276] <= 32'd3352;
		word[15'd4277] <= 32'd3353;
		word[15'd4278] <= 32'd3354;
		word[15'd4279] <= 32'd3355;
		word[15'd4280] <= 32'd3356;
		word[15'd4281] <= 32'd3357;
		word[15'd4282] <= 32'd3358;
		word[15'd4283] <= 32'd3359;
		word[15'd4284] <= 32'd3360;
		word[15'd4285] <= 32'd3361;
		word[15'd4286] <= 32'd3362;
		word[15'd4287] <= 32'd3363;
		word[15'd4288] <= 32'd3364;
		word[15'd4289] <= 32'd3365;
		word[15'd4290] <= 32'd3366;
		word[15'd4291] <= 32'd3367;
		word[15'd4292] <= 32'd3368;
		word[15'd4293] <= 32'd3369;
		word[15'd4294] <= 32'd3370;
		word[15'd4295] <= 32'd3371;
		word[15'd4296] <= 32'd3372;
		word[15'd4297] <= 32'd3373;
		word[15'd4298] <= 32'd3374;
		word[15'd4299] <= 32'd3375;
		word[15'd4300] <= 32'd3376;
		word[15'd4301] <= 32'd3377;
		word[15'd4302] <= 32'd3378;
		word[15'd4303] <= 32'd3379;
		word[15'd4304] <= 32'd3380;
		word[15'd4305] <= 32'd3381;
		word[15'd4306] <= 32'd3382;
		word[15'd4307] <= 32'd3383;
		word[15'd4308] <= 32'd3384;
		word[15'd4309] <= 32'd3385;
		word[15'd4310] <= 32'd3386;
		word[15'd4311] <= 32'd3387;
		word[15'd4312] <= 32'd3388;
		word[15'd4313] <= 32'd3389;
		word[15'd4314] <= 32'd3390;
		word[15'd4315] <= 32'd3391;
		word[15'd4316] <= 32'd3392;
		word[15'd4317] <= 32'd3393;
		word[15'd4318] <= 32'd3394;
		word[15'd4319] <= 32'd3395;
		word[15'd4320] <= 32'd3396;
		word[15'd4321] <= 32'd3397;
		word[15'd4322] <= 32'd3398;
		word[15'd4323] <= 32'd3399;
		word[15'd4324] <= 32'd3400;
		word[15'd4325] <= 32'd3401;
		word[15'd4326] <= 32'd3402;
		word[15'd4327] <= 32'd3403;
		word[15'd4328] <= 32'd3404;
		word[15'd4329] <= 32'd3405;
		word[15'd4330] <= 32'd3406;
		word[15'd4331] <= 32'd3407;
		word[15'd4332] <= 32'd3408;
		word[15'd4333] <= 32'd3409;
		word[15'd4334] <= 32'd3410;
		word[15'd4335] <= 32'd3411;
		word[15'd4336] <= 32'd3412;
		word[15'd4337] <= 32'd3413;
		word[15'd4338] <= 32'd3414;
		word[15'd4339] <= 32'd3415;
		word[15'd4340] <= 32'd3416;
		word[15'd4341] <= 32'd3417;
		word[15'd4342] <= 32'd3418;
		word[15'd4343] <= 32'd3419;
		word[15'd4344] <= 32'd3420;
		word[15'd4345] <= 32'd3421;
		word[15'd4346] <= 32'd3422;
		word[15'd4347] <= 32'd3423;
		word[15'd4348] <= 32'd3424;
		word[15'd4349] <= 32'd3425;
		word[15'd4350] <= 32'd3426;
		word[15'd4351] <= 32'd3427;
		word[15'd4352] <= 32'd3428;
		word[15'd4353] <= 32'd3429;
		word[15'd4354] <= 32'd3430;
		word[15'd4355] <= 32'd3431;
		word[15'd4356] <= 32'd3432;
		word[15'd4357] <= 32'd3433;
		word[15'd4358] <= 32'd3434;
		word[15'd4359] <= 32'd3435;
		word[15'd4360] <= 32'd3436;
		word[15'd4361] <= 32'd3437;
		word[15'd4362] <= 32'd3438;
		word[15'd4363] <= 32'd3439;
		word[15'd4364] <= 32'd3440;
		word[15'd4365] <= 32'd3441;
		word[15'd4366] <= 32'd3442;
		word[15'd4367] <= 32'd3443;
		word[15'd4368] <= 32'd3444;
		word[15'd4369] <= 32'd3445;
		word[15'd4370] <= 32'd3446;
		word[15'd4371] <= 32'd3447;
		word[15'd4372] <= 32'd3448;
		word[15'd4373] <= 32'd3449;
		word[15'd4374] <= 32'd3450;
		word[15'd4375] <= 32'd3451;
		word[15'd4376] <= 32'd3452;
		word[15'd4377] <= 32'd3453;
		word[15'd4378] <= 32'd3454;
		word[15'd4379] <= 32'd3455;
		word[15'd4380] <= 32'd3456;
		word[15'd4381] <= 32'd3457;
		word[15'd4382] <= 32'd3458;
		word[15'd4383] <= 32'd3459;
		word[15'd4384] <= 32'd3460;
		word[15'd4385] <= 32'd3461;
		word[15'd4386] <= 32'd3462;
		word[15'd4387] <= 32'd3463;
		word[15'd4388] <= 32'd3464;
		word[15'd4389] <= 32'd3465;
		word[15'd4390] <= 32'd3466;
		word[15'd4391] <= 32'd3467;
		word[15'd4392] <= 32'd3468;
		word[15'd4393] <= 32'd3469;
		word[15'd4394] <= 32'd3470;
		word[15'd4395] <= 32'd3471;
		word[15'd4396] <= 32'd3472;
		word[15'd4397] <= 32'd3473;
		word[15'd4398] <= 32'd3474;
		word[15'd4399] <= 32'd3475;
		word[15'd4400] <= 32'd3476;
		word[15'd4401] <= 32'd3477;
		word[15'd4402] <= 32'd3478;
		word[15'd4403] <= 32'd3479;
		word[15'd4404] <= 32'd3480;
		word[15'd4405] <= 32'd3481;
		word[15'd4406] <= 32'd3482;
		word[15'd4407] <= 32'd3483;
		word[15'd4408] <= 32'd3484;
		word[15'd4409] <= 32'd3485;
		word[15'd4410] <= 32'd3486;
		word[15'd4411] <= 32'd3487;
		word[15'd4412] <= 32'd3488;
		word[15'd4413] <= 32'd3489;
		word[15'd4414] <= 32'd3490;
		word[15'd4415] <= 32'd3491;
		word[15'd4416] <= 32'd3492;
		word[15'd4417] <= 32'd3493;
		word[15'd4418] <= 32'd3494;
		word[15'd4419] <= 32'd3495;
		word[15'd4420] <= 32'd3496;
		word[15'd4421] <= 32'd3497;
		word[15'd4422] <= 32'd3498;
		word[15'd4423] <= 32'd3499;
		word[15'd4424] <= 32'd3500;
		word[15'd4425] <= 32'd3501;
		word[15'd4426] <= 32'd3502;
		word[15'd4427] <= 32'd3503;
		word[15'd4428] <= 32'd3504;
		word[15'd4429] <= 32'd3505;
		word[15'd4430] <= 32'd3506;
		word[15'd4431] <= 32'd3507;
		word[15'd4432] <= 32'd3508;
		word[15'd4433] <= 32'd3509;
		word[15'd4434] <= 32'd3510;
		word[15'd4435] <= 32'd3511;
		word[15'd4436] <= 32'd3512;
		word[15'd4437] <= 32'd3513;
		word[15'd4438] <= 32'd3514;
		word[15'd4439] <= 32'd3515;
		word[15'd4440] <= 32'd3516;
		word[15'd4441] <= 32'd3517;
		word[15'd4442] <= 32'd3518;
		word[15'd4443] <= 32'd3519;
		word[15'd4444] <= 32'd3520;
		word[15'd4445] <= 32'd3521;
		word[15'd4446] <= 32'd3522;
		word[15'd4447] <= 32'd3523;
		word[15'd4448] <= 32'd3524;
		word[15'd4449] <= 32'd3525;
		word[15'd4450] <= 32'd3526;
		word[15'd4451] <= 32'd3527;
		word[15'd4452] <= 32'd3528;
		word[15'd4453] <= 32'd3529;
		word[15'd4454] <= 32'd3530;
		word[15'd4455] <= 32'd3531;
		word[15'd4456] <= 32'd3532;
		word[15'd4457] <= 32'd3533;
		word[15'd4458] <= 32'd3534;
		word[15'd4459] <= 32'd3535;
		word[15'd4460] <= 32'd3536;
		word[15'd4461] <= 32'd3537;
		word[15'd4462] <= 32'd3538;
		word[15'd4463] <= 32'd3539;
		word[15'd4464] <= 32'd3540;
		word[15'd4465] <= 32'd3541;
		word[15'd4466] <= 32'd3542;
		word[15'd4467] <= 32'd3543;
		word[15'd4468] <= 32'd3544;
		word[15'd4469] <= 32'd3545;
		word[15'd4470] <= 32'd3546;
		word[15'd4471] <= 32'd3547;
		word[15'd4472] <= 32'd3548;
		word[15'd4473] <= 32'd3549;
		word[15'd4474] <= 32'd3550;
		word[15'd4475] <= 32'd3551;
		word[15'd4476] <= 32'd3552;
		word[15'd4477] <= 32'd3553;
		word[15'd4478] <= 32'd3554;
		word[15'd4479] <= 32'd3555;
		word[15'd4480] <= 32'd3556;
		word[15'd4481] <= 32'd3557;
		word[15'd4482] <= 32'd3558;
		word[15'd4483] <= 32'd3559;
		word[15'd4484] <= 32'd3560;
		word[15'd4485] <= 32'd3561;
		word[15'd4486] <= 32'd3562;
		word[15'd4487] <= 32'd3563;
		word[15'd4488] <= 32'd3564;
		word[15'd4489] <= 32'd3565;
		word[15'd4490] <= 32'd3566;
		word[15'd4491] <= 32'd3567;
		word[15'd4492] <= 32'd3568;
		word[15'd4493] <= 32'd3569;
		word[15'd4494] <= 32'd3570;
		word[15'd4495] <= 32'd3571;
		word[15'd4496] <= 32'd3572;
		word[15'd4497] <= 32'd3573;
		word[15'd4498] <= 32'd3574;
		word[15'd4499] <= 32'd3575;
		word[15'd4500] <= 32'd3576;
		word[15'd4501] <= 32'd3577;
		word[15'd4502] <= 32'd3578;
		word[15'd4503] <= 32'd3579;
		word[15'd4504] <= 32'd3580;
		word[15'd4505] <= 32'd3581;
		word[15'd4506] <= 32'd3582;
		word[15'd4507] <= 32'd3583;
		word[15'd4508] <= 32'd3584;
		word[15'd4509] <= 32'd3585;
		word[15'd4510] <= 32'd3586;
		word[15'd4511] <= 32'd3587;
		word[15'd4512] <= 32'd3588;
		word[15'd4513] <= 32'd3589;
		word[15'd4514] <= 32'd3590;
		word[15'd4515] <= 32'd3591;
		word[15'd4516] <= 32'd3592;
		word[15'd4517] <= 32'd3593;
		word[15'd4518] <= 32'd3594;
		word[15'd4519] <= 32'd3595;
		word[15'd4520] <= 32'd3596;
		word[15'd4521] <= 32'd3597;
		word[15'd4522] <= 32'd3598;
		word[15'd4523] <= 32'd3599;
		word[15'd4524] <= 32'd3600;
		word[15'd4525] <= 32'd3601;
		word[15'd4526] <= 32'd3602;
		word[15'd4527] <= 32'd3603;
		word[15'd4528] <= 32'd3604;
		word[15'd4529] <= 32'd3605;
		word[15'd4530] <= 32'd3606;
		word[15'd4531] <= 32'd3607;
		word[15'd4532] <= 32'd3608;
		word[15'd4533] <= 32'd3609;
		word[15'd4534] <= 32'd3610;
		word[15'd4535] <= 32'd3611;
		word[15'd4536] <= 32'd3612;
		word[15'd4537] <= 32'd3613;
		word[15'd4538] <= 32'd3614;
		word[15'd4539] <= 32'd3615;
		word[15'd4540] <= 32'd3616;
		word[15'd4541] <= 32'd3617;
		word[15'd4542] <= 32'd3618;
		word[15'd4543] <= 32'd3619;
		word[15'd4544] <= 32'd3620;
		word[15'd4545] <= 32'd3621;
		word[15'd4546] <= 32'd3622;
		word[15'd4547] <= 32'd3623;
		word[15'd4548] <= 32'd3624;
		word[15'd4549] <= 32'd3625;
		word[15'd4550] <= 32'd3626;
		word[15'd4551] <= 32'd3627;
		word[15'd4552] <= 32'd3628;
		word[15'd4553] <= 32'd3629;
		word[15'd4554] <= 32'd3630;
		word[15'd4555] <= 32'd3631;
		word[15'd4556] <= 32'd3632;
		word[15'd4557] <= 32'd3633;
		word[15'd4558] <= 32'd3634;
		word[15'd4559] <= 32'd3635;
		word[15'd4560] <= 32'd3636;
		word[15'd4561] <= 32'd3637;
		word[15'd4562] <= 32'd3638;
		word[15'd4563] <= 32'd3639;
		word[15'd4564] <= 32'd3640;
		word[15'd4565] <= 32'd3641;
		word[15'd4566] <= 32'd3642;
		word[15'd4567] <= 32'd3643;
		word[15'd4568] <= 32'd3644;
		word[15'd4569] <= 32'd3645;
		word[15'd4570] <= 32'd3646;
		word[15'd4571] <= 32'd3647;
		word[15'd4572] <= 32'd3648;
		word[15'd4573] <= 32'd3649;
		word[15'd4574] <= 32'd3650;
		word[15'd4575] <= 32'd3651;
		word[15'd4576] <= 32'd3652;
		word[15'd4577] <= 32'd3653;
		word[15'd4578] <= 32'd3654;
		word[15'd4579] <= 32'd3655;
		word[15'd4580] <= 32'd3656;
		word[15'd4581] <= 32'd3657;
		word[15'd4582] <= 32'd3658;
		word[15'd4583] <= 32'd3659;
		word[15'd4584] <= 32'd3660;
		word[15'd4585] <= 32'd3661;
		word[15'd4586] <= 32'd3662;
		word[15'd4587] <= 32'd3663;
		word[15'd4588] <= 32'd3664;
		word[15'd4589] <= 32'd3665;
		word[15'd4590] <= 32'd3666;
		word[15'd4591] <= 32'd3667;
		word[15'd4592] <= 32'd3668;
		word[15'd4593] <= 32'd3669;
		word[15'd4594] <= 32'd3670;
		word[15'd4595] <= 32'd3671;
		word[15'd4596] <= 32'd3672;
		word[15'd4597] <= 32'd3673;
		word[15'd4598] <= 32'd3674;
		word[15'd4599] <= 32'd3675;
		word[15'd4600] <= 32'd3676;
		word[15'd4601] <= 32'd3677;
		word[15'd4602] <= 32'd3678;
		word[15'd4603] <= 32'd3679;
		word[15'd4604] <= 32'd3680;
		word[15'd4605] <= 32'd3681;
		word[15'd4606] <= 32'd3682;
		word[15'd4607] <= 32'd3683;
		word[15'd4608] <= 32'd3684;
		word[15'd4609] <= 32'd3685;
		word[15'd4610] <= 32'd3686;
		word[15'd4611] <= 32'd3687;
		word[15'd4612] <= 32'd3688;
		word[15'd4613] <= 32'd3689;
		word[15'd4614] <= 32'd3690;
		word[15'd4615] <= 32'd3691;
		word[15'd4616] <= 32'd3692;
		word[15'd4617] <= 32'd3693;
		word[15'd4618] <= 32'd3694;
		word[15'd4619] <= 32'd3695;
		word[15'd4620] <= 32'd3696;
		word[15'd4621] <= 32'd3697;
		word[15'd4622] <= 32'd3698;
		word[15'd4623] <= 32'd3699;
		word[15'd4624] <= 32'd3700;
		word[15'd4625] <= 32'd3701;
		word[15'd4626] <= 32'd3702;
		word[15'd4627] <= 32'd3703;
		word[15'd4628] <= 32'd3704;
		word[15'd4629] <= 32'd3705;
		word[15'd4630] <= 32'd3706;
		word[15'd4631] <= 32'd3707;
		word[15'd4632] <= 32'd3708;
		word[15'd4633] <= 32'd3709;
		word[15'd4634] <= 32'd3710;
		word[15'd4635] <= 32'd3711;
		word[15'd4636] <= 32'd3712;
		word[15'd4637] <= 32'd3713;
		word[15'd4638] <= 32'd3714;
		word[15'd4639] <= 32'd3715;
		word[15'd4640] <= 32'd3716;
		word[15'd4641] <= 32'd3717;
		word[15'd4642] <= 32'd3718;
		word[15'd4643] <= 32'd3719;
		word[15'd4644] <= 32'd3720;
		word[15'd4645] <= 32'd3721;
		word[15'd4646] <= 32'd3722;
		word[15'd4647] <= 32'd3723;
		word[15'd4648] <= 32'd3724;
		word[15'd4649] <= 32'd3725;
		word[15'd4650] <= 32'd3726;
		word[15'd4651] <= 32'd3727;
		word[15'd4652] <= 32'd3728;
		word[15'd4653] <= 32'd3729;
		word[15'd4654] <= 32'd3730;
		word[15'd4655] <= 32'd3731;
		word[15'd4656] <= 32'd3732;
		word[15'd4657] <= 32'd3733;
		word[15'd4658] <= 32'd3734;
		word[15'd4659] <= 32'd3735;
		word[15'd4660] <= 32'd3736;
		word[15'd4661] <= 32'd3737;
		word[15'd4662] <= 32'd3738;
		word[15'd4663] <= 32'd3739;
		word[15'd4664] <= 32'd3740;
		word[15'd4665] <= 32'd3741;
		word[15'd4666] <= 32'd3742;
		word[15'd4667] <= 32'd3743;
		word[15'd4668] <= 32'd3744;
		word[15'd4669] <= 32'd3745;
		word[15'd4670] <= 32'd3746;
		word[15'd4671] <= 32'd3747;
		word[15'd4672] <= 32'd3748;
		word[15'd4673] <= 32'd3749;
		word[15'd4674] <= 32'd3750;
		word[15'd4675] <= 32'd3751;
		word[15'd4676] <= 32'd3752;
		word[15'd4677] <= 32'd3753;
		word[15'd4678] <= 32'd3754;
		word[15'd4679] <= 32'd3755;
		word[15'd4680] <= 32'd3756;
		word[15'd4681] <= 32'd3757;
		word[15'd4682] <= 32'd3758;
		word[15'd4683] <= 32'd3759;
		word[15'd4684] <= 32'd3760;
		word[15'd4685] <= 32'd3761;
		word[15'd4686] <= 32'd3762;
		word[15'd4687] <= 32'd3763;
		word[15'd4688] <= 32'd3764;
		word[15'd4689] <= 32'd3765;
		word[15'd4690] <= 32'd3766;
		word[15'd4691] <= 32'd3767;
		word[15'd4692] <= 32'd3768;
		word[15'd4693] <= 32'd3769;
		word[15'd4694] <= 32'd3770;
		word[15'd4695] <= 32'd3771;
		word[15'd4696] <= 32'd3772;
		word[15'd4697] <= 32'd3773;
		word[15'd4698] <= 32'd3774;
		word[15'd4699] <= 32'd3775;
		word[15'd4700] <= 32'd3776;
		word[15'd4701] <= 32'd3777;
		word[15'd4702] <= 32'd3778;
		word[15'd4703] <= 32'd3779;
		word[15'd4704] <= 32'd3780;
		word[15'd4705] <= 32'd3781;
		word[15'd4706] <= 32'd3782;
		word[15'd4707] <= 32'd3783;
		word[15'd4708] <= 32'd3784;
		word[15'd4709] <= 32'd3785;
		word[15'd4710] <= 32'd3786;
		word[15'd4711] <= 32'd3787;
		word[15'd4712] <= 32'd3788;
		word[15'd4713] <= 32'd3789;
		word[15'd4714] <= 32'd3790;
		word[15'd4715] <= 32'd3791;
		word[15'd4716] <= 32'd3792;
		word[15'd4717] <= 32'd3793;
		word[15'd4718] <= 32'd3794;
		word[15'd4719] <= 32'd3795;
		word[15'd4720] <= 32'd3796;
		word[15'd4721] <= 32'd3797;
		word[15'd4722] <= 32'd3798;
		word[15'd4723] <= 32'd3799;
		word[15'd4724] <= 32'd3800;
		word[15'd4725] <= 32'd3801;
		word[15'd4726] <= 32'd3802;
		word[15'd4727] <= 32'd3803;
		word[15'd4728] <= 32'd3804;
		word[15'd4729] <= 32'd3805;
		word[15'd4730] <= 32'd3806;
		word[15'd4731] <= 32'd3807;
		word[15'd4732] <= 32'd3808;
		word[15'd4733] <= 32'd3809;
		word[15'd4734] <= 32'd3810;
		word[15'd4735] <= 32'd3811;
		word[15'd4736] <= 32'd3812;
		word[15'd4737] <= 32'd3813;
		word[15'd4738] <= 32'd3814;
		word[15'd4739] <= 32'd3815;
		word[15'd4740] <= 32'd3816;
		word[15'd4741] <= 32'd3817;
		word[15'd4742] <= 32'd3818;
		word[15'd4743] <= 32'd3819;
		word[15'd4744] <= 32'd3820;
		word[15'd4745] <= 32'd3821;
		word[15'd4746] <= 32'd3822;
		word[15'd4747] <= 32'd3823;
		word[15'd4748] <= 32'd3824;
		word[15'd4749] <= 32'd3825;
		word[15'd4750] <= 32'd3826;
		word[15'd4751] <= 32'd3827;
		word[15'd4752] <= 32'd3828;
		word[15'd4753] <= 32'd3829;
		word[15'd4754] <= 32'd3830;
		word[15'd4755] <= 32'd3831;
		word[15'd4756] <= 32'd3832;
		word[15'd4757] <= 32'd3833;
		word[15'd4758] <= 32'd3834;
		word[15'd4759] <= 32'd3835;
		word[15'd4760] <= 32'd3836;
		word[15'd4761] <= 32'd3837;
		word[15'd4762] <= 32'd3838;
		word[15'd4763] <= 32'd3839;
		word[15'd4764] <= 32'd3840;
		word[15'd4765] <= 32'd3841;
		word[15'd4766] <= 32'd3842;
		word[15'd4767] <= 32'd3843;
		word[15'd4768] <= 32'd3844;
		word[15'd4769] <= 32'd3845;
		word[15'd4770] <= 32'd3846;
		word[15'd4771] <= 32'd3847;
		word[15'd4772] <= 32'd3848;
		word[15'd4773] <= 32'd3849;
		word[15'd4774] <= 32'd3850;
		word[15'd4775] <= 32'd3851;
		word[15'd4776] <= 32'd3852;
		word[15'd4777] <= 32'd3853;
		word[15'd4778] <= 32'd3854;
		word[15'd4779] <= 32'd3855;
		word[15'd4780] <= 32'd3856;
		word[15'd4781] <= 32'd3857;
		word[15'd4782] <= 32'd3858;
		word[15'd4783] <= 32'd3859;
		word[15'd4784] <= 32'd3860;
		word[15'd4785] <= 32'd3861;
		word[15'd4786] <= 32'd3862;
		word[15'd4787] <= 32'd3863;
		word[15'd4788] <= 32'd3864;
		word[15'd4789] <= 32'd3865;
		word[15'd4790] <= 32'd3866;
		word[15'd4791] <= 32'd3867;
		word[15'd4792] <= 32'd3868;
		word[15'd4793] <= 32'd3869;
		word[15'd4794] <= 32'd3870;
		word[15'd4795] <= 32'd3871;
		word[15'd4796] <= 32'd3872;
		word[15'd4797] <= 32'd3873;
		word[15'd4798] <= 32'd3874;
		word[15'd4799] <= 32'd3875;
		word[15'd4800] <= 32'd3876;
		word[15'd4801] <= 32'd3877;
		word[15'd4802] <= 32'd3878;
		word[15'd4803] <= 32'd3879;
		word[15'd4804] <= 32'd3880;
		word[15'd4805] <= 32'd3881;
		word[15'd4806] <= 32'd3882;
		word[15'd4807] <= 32'd3883;
		word[15'd4808] <= 32'd3884;
		word[15'd4809] <= 32'd3885;
		word[15'd4810] <= 32'd3886;
		word[15'd4811] <= 32'd3887;
		word[15'd4812] <= 32'd3888;
		word[15'd4813] <= 32'd3889;
		word[15'd4814] <= 32'd3890;
		word[15'd4815] <= 32'd3891;
		word[15'd4816] <= 32'd3892;
		word[15'd4817] <= 32'd3893;
		word[15'd4818] <= 32'd3894;
		word[15'd4819] <= 32'd3895;
		word[15'd4820] <= 32'd3896;
		word[15'd4821] <= 32'd3897;
		word[15'd4822] <= 32'd3898;
		word[15'd4823] <= 32'd3899;
		word[15'd4824] <= 32'd3900;
		word[15'd4825] <= 32'd3901;
		word[15'd4826] <= 32'd3902;
		word[15'd4827] <= 32'd3903;
		word[15'd4828] <= 32'd3904;
		word[15'd4829] <= 32'd3905;
		word[15'd4830] <= 32'd3906;
		word[15'd4831] <= 32'd3907;
		word[15'd4832] <= 32'd3908;
		word[15'd4833] <= 32'd3909;
		word[15'd4834] <= 32'd3910;
		word[15'd4835] <= 32'd3911;
		word[15'd4836] <= 32'd3912;
		word[15'd4837] <= 32'd3913;
		word[15'd4838] <= 32'd3914;
		word[15'd4839] <= 32'd3915;
		word[15'd4840] <= 32'd3916;
		word[15'd4841] <= 32'd3917;
		word[15'd4842] <= 32'd3918;
		word[15'd4843] <= 32'd3919;
		word[15'd4844] <= 32'd3920;
		word[15'd4845] <= 32'd3921;
		word[15'd4846] <= 32'd3922;
		word[15'd4847] <= 32'd3923;
		word[15'd4848] <= 32'd3924;
		word[15'd4849] <= 32'd3925;
		word[15'd4850] <= 32'd3926;
		word[15'd4851] <= 32'd3927;
		word[15'd4852] <= 32'd3928;
		word[15'd4853] <= 32'd3929;
		word[15'd4854] <= 32'd3930;
		word[15'd4855] <= 32'd3931;
		word[15'd4856] <= 32'd3932;
		word[15'd4857] <= 32'd3933;
		word[15'd4858] <= 32'd3934;
		word[15'd4859] <= 32'd3935;
		word[15'd4860] <= 32'd3936;
		word[15'd4861] <= 32'd3937;
		word[15'd4862] <= 32'd3938;
		word[15'd4863] <= 32'd3939;
		word[15'd4864] <= 32'd3940;
		word[15'd4865] <= 32'd3941;
		word[15'd4866] <= 32'd3942;
		word[15'd4867] <= 32'd3943;
		word[15'd4868] <= 32'd3944;
		word[15'd4869] <= 32'd3945;
		word[15'd4870] <= 32'd3946;
		word[15'd4871] <= 32'd3947;
		word[15'd4872] <= 32'd3948;
		word[15'd4873] <= 32'd3949;
		word[15'd4874] <= 32'd3950;
		word[15'd4875] <= 32'd3951;
		word[15'd4876] <= 32'd3952;
		word[15'd4877] <= 32'd3953;
		word[15'd4878] <= 32'd3954;
		word[15'd4879] <= 32'd3955;
		word[15'd4880] <= 32'd3956;
		word[15'd4881] <= 32'd3957;
		word[15'd4882] <= 32'd3958;
		word[15'd4883] <= 32'd3959;
		word[15'd4884] <= 32'd3960;
		word[15'd4885] <= 32'd3961;
		word[15'd4886] <= 32'd3962;
		word[15'd4887] <= 32'd3963;
		word[15'd4888] <= 32'd3964;
		word[15'd4889] <= 32'd3965;
		word[15'd4890] <= 32'd3966;
		word[15'd4891] <= 32'd3967;
		word[15'd4892] <= 32'd3968;
		word[15'd4893] <= 32'd3969;
		word[15'd4894] <= 32'd3970;
		word[15'd4895] <= 32'd3971;
		word[15'd4896] <= 32'd3972;
		word[15'd4897] <= 32'd3973;
		word[15'd4898] <= 32'd3974;
		word[15'd4899] <= 32'd3975;
		word[15'd4900] <= 32'd3976;
		word[15'd4901] <= 32'd3977;
		word[15'd4902] <= 32'd3978;
		word[15'd4903] <= 32'd3979;
		word[15'd4904] <= 32'd3980;
		word[15'd4905] <= 32'd3981;
		word[15'd4906] <= 32'd3982;
		word[15'd4907] <= 32'd3983;
		word[15'd4908] <= 32'd3984;
		word[15'd4909] <= 32'd3985;
		word[15'd4910] <= 32'd3986;
		word[15'd4911] <= 32'd3987;
		word[15'd4912] <= 32'd3988;
		word[15'd4913] <= 32'd3989;
		word[15'd4914] <= 32'd3990;
		word[15'd4915] <= 32'd3991;
		word[15'd4916] <= 32'd3992;
		word[15'd4917] <= 32'd3993;
		word[15'd4918] <= 32'd3994;
		word[15'd4919] <= 32'd3995;
		word[15'd4920] <= 32'd3996;
		word[15'd4921] <= 32'd3997;
		word[15'd4922] <= 32'd3998;
		word[15'd4923] <= 32'd3999;
		word[15'd4924] <= 32'd4000;
		word[15'd4925] <= 32'd4001;
		word[15'd4926] <= 32'd4002;
		word[15'd4927] <= 32'd4003;
		word[15'd4928] <= 32'd4004;
		word[15'd4929] <= 32'd4005;
		word[15'd4930] <= 32'd4006;
		word[15'd4931] <= 32'd4007;
		word[15'd4932] <= 32'd4008;
		word[15'd4933] <= 32'd4009;
		word[15'd4934] <= 32'd4010;
		word[15'd4935] <= 32'd4011;
		word[15'd4936] <= 32'd4012;
		word[15'd4937] <= 32'd4013;
		word[15'd4938] <= 32'd4014;
		word[15'd4939] <= 32'd4015;
		word[15'd4940] <= 32'd4016;
		word[15'd4941] <= 32'd4017;
		word[15'd4942] <= 32'd4018;
		word[15'd4943] <= 32'd4019;
		word[15'd4944] <= 32'd4020;
		word[15'd4945] <= 32'd4021;
		word[15'd4946] <= 32'd4022;
		word[15'd4947] <= 32'd4023;
		word[15'd4948] <= 32'd4024;
		word[15'd4949] <= 32'd4025;
		word[15'd4950] <= 32'd4026;
		word[15'd4951] <= 32'd4027;
		word[15'd4952] <= 32'd4028;
		word[15'd4953] <= 32'd4029;
		word[15'd4954] <= 32'd4030;
		word[15'd4955] <= 32'd4031;
		word[15'd4956] <= 32'd4032;
		word[15'd4957] <= 32'd4033;
		word[15'd4958] <= 32'd4034;
		word[15'd4959] <= 32'd4035;
		word[15'd4960] <= 32'd4036;
		word[15'd4961] <= 32'd4037;
		word[15'd4962] <= 32'd4038;
		word[15'd4963] <= 32'd4039;
		word[15'd4964] <= 32'd4040;
		word[15'd4965] <= 32'd4041;
		word[15'd4966] <= 32'd4042;
		word[15'd4967] <= 32'd4043;
		word[15'd4968] <= 32'd4044;
		word[15'd4969] <= 32'd4045;
		word[15'd4970] <= 32'd4046;
		word[15'd4971] <= 32'd4047;
		word[15'd4972] <= 32'd4048;
		word[15'd4973] <= 32'd4049;
		word[15'd4974] <= 32'd4050;
		word[15'd4975] <= 32'd4051;
		word[15'd4976] <= 32'd4052;
		word[15'd4977] <= 32'd4053;
		word[15'd4978] <= 32'd4054;
		word[15'd4979] <= 32'd4055;
		word[15'd4980] <= 32'd4056;
		word[15'd4981] <= 32'd4057;
		word[15'd4982] <= 32'd4058;
		word[15'd4983] <= 32'd4059;
		word[15'd4984] <= 32'd4060;
		word[15'd4985] <= 32'd4061;
		word[15'd4986] <= 32'd4062;
		word[15'd4987] <= 32'd4063;
		word[15'd4988] <= 32'd4064;
		word[15'd4989] <= 32'd4065;
		word[15'd4990] <= 32'd4066;
		word[15'd4991] <= 32'd4067;
		word[15'd4992] <= 32'd4068;
		word[15'd4993] <= 32'd4069;
		word[15'd4994] <= 32'd4070;
		word[15'd4995] <= 32'd4071;
		word[15'd4996] <= 32'd4072;
		word[15'd4997] <= 32'd4073;
		word[15'd4998] <= 32'd4074;
		word[15'd4999] <= 32'd4075;
		word[15'd5000] <= 32'd4076;
		word[15'd5001] <= 32'd4077;
		word[15'd5002] <= 32'd4078;
		word[15'd5003] <= 32'd4079;
		word[15'd5004] <= 32'd4080;
		word[15'd5005] <= 32'd4081;
		word[15'd5006] <= 32'd4082;
		word[15'd5007] <= 32'd4083;
		word[15'd5008] <= 32'd4084;
		word[15'd5009] <= 32'd4085;
		word[15'd5010] <= 32'd4086;
		word[15'd5011] <= 32'd4087;
		word[15'd5012] <= 32'd4088;
		word[15'd5013] <= 32'd4089;
		word[15'd5014] <= 32'd4090;
		word[15'd5015] <= 32'd4091;
		word[15'd5016] <= 32'd4092;
		word[15'd5017] <= 32'd4093;
		word[15'd5018] <= 32'd4094;
		word[15'd5019] <= 32'd4095;
		word[15'd5020] <= 32'd4096;
		word[15'd5021] <= 32'd4097;
		word[15'd5022] <= 32'd4098;
		word[15'd5023] <= 32'd4099;
		word[15'd5024] <= 32'd4100;
		word[15'd5025] <= 32'd4101;
		word[15'd5026] <= 32'd4102;
		word[15'd5027] <= 32'd4103;
		word[15'd5028] <= 32'd4104;
		word[15'd5029] <= 32'd4105;
		word[15'd5030] <= 32'd4106;
		word[15'd5031] <= 32'd4107;
		word[15'd5032] <= 32'd4108;
		word[15'd5033] <= 32'd4109;
		word[15'd5034] <= 32'd4110;
		word[15'd5035] <= 32'd4111;
		word[15'd5036] <= 32'd4112;
		word[15'd5037] <= 32'd4113;
		word[15'd5038] <= 32'd4114;
		word[15'd5039] <= 32'd4115;
		word[15'd5040] <= 32'd4116;
		word[15'd5041] <= 32'd4117;
		word[15'd5042] <= 32'd4118;
		word[15'd5043] <= 32'd4119;
		word[15'd5044] <= 32'd4120;
		word[15'd5045] <= 32'd4121;
		word[15'd5046] <= 32'd4122;
		word[15'd5047] <= 32'd4123;
		word[15'd5048] <= 32'd4124;
		word[15'd5049] <= 32'd4125;
		word[15'd5050] <= 32'd4126;
		word[15'd5051] <= 32'd4127;
		word[15'd5052] <= 32'd4128;
		word[15'd5053] <= 32'd4129;
		word[15'd5054] <= 32'd4130;
		word[15'd5055] <= 32'd4131;
		word[15'd5056] <= 32'd4132;
		word[15'd5057] <= 32'd4133;
		word[15'd5058] <= 32'd4134;
		word[15'd5059] <= 32'd4135;
		word[15'd5060] <= 32'd4136;
		word[15'd5061] <= 32'd4137;
		word[15'd5062] <= 32'd4138;
		word[15'd5063] <= 32'd4139;
		word[15'd5064] <= 32'd4140;
		word[15'd5065] <= 32'd4141;
		word[15'd5066] <= 32'd4142;
		word[15'd5067] <= 32'd4143;
		word[15'd5068] <= 32'd4144;
		word[15'd5069] <= 32'd4145;
		word[15'd5070] <= 32'd4146;
		word[15'd5071] <= 32'd4147;
		word[15'd5072] <= 32'd4148;
		word[15'd5073] <= 32'd4149;
		word[15'd5074] <= 32'd4150;
		word[15'd5075] <= 32'd4151;
		word[15'd5076] <= 32'd4152;
		word[15'd5077] <= 32'd4153;
		word[15'd5078] <= 32'd4154;
		word[15'd5079] <= 32'd4155;
		word[15'd5080] <= 32'd4156;
		word[15'd5081] <= 32'd4157;
		word[15'd5082] <= 32'd4158;
		word[15'd5083] <= 32'd4159;
		word[15'd5084] <= 32'd4160;
		word[15'd5085] <= 32'd4161;
		word[15'd5086] <= 32'd4162;
		word[15'd5087] <= 32'd4163;
		word[15'd5088] <= 32'd4164;
		word[15'd5089] <= 32'd4165;
		word[15'd5090] <= 32'd4166;
		word[15'd5091] <= 32'd4167;
		word[15'd5092] <= 32'd4168;
		word[15'd5093] <= 32'd4169;
		word[15'd5094] <= 32'd4170;
		word[15'd5095] <= 32'd4171;
		word[15'd5096] <= 32'd4172;
		word[15'd5097] <= 32'd4173;
		word[15'd5098] <= 32'd4174;
		word[15'd5099] <= 32'd4175;
		word[15'd5100] <= 32'd4176;
		word[15'd5101] <= 32'd4177;
		word[15'd5102] <= 32'd4178;
		word[15'd5103] <= 32'd4179;
		word[15'd5104] <= 32'd4180;
		word[15'd5105] <= 32'd4181;
		word[15'd5106] <= 32'd4182;
		word[15'd5107] <= 32'd4183;
		word[15'd5108] <= 32'd4184;
		word[15'd5109] <= 32'd4185;
		word[15'd5110] <= 32'd4186;
		word[15'd5111] <= 32'd4187;
		word[15'd5112] <= 32'd4188;
		word[15'd5113] <= 32'd4189;
		word[15'd5114] <= 32'd4190;
		word[15'd5115] <= 32'd4191;
		word[15'd5116] <= 32'd4192;
		word[15'd5117] <= 32'd4193;
		word[15'd5118] <= 32'd4194;
		word[15'd5119] <= 32'd4195;
		word[15'd5120] <= 32'd4196;
		word[15'd5121] <= 32'd4197;
		word[15'd5122] <= 32'd4198;
		word[15'd5123] <= 32'd4199;
		word[15'd5124] <= 32'd4200;
		word[15'd5125] <= 32'd4201;
		word[15'd5126] <= 32'd4202;
		word[15'd5127] <= 32'd4203;
		word[15'd5128] <= 32'd4204;
		word[15'd5129] <= 32'd4205;
		word[15'd5130] <= 32'd4206;
		word[15'd5131] <= 32'd4207;
		word[15'd5132] <= 32'd4208;
		word[15'd5133] <= 32'd4209;
		word[15'd5134] <= 32'd4210;
		word[15'd5135] <= 32'd4211;
		word[15'd5136] <= 32'd4212;
		word[15'd5137] <= 32'd4213;
		word[15'd5138] <= 32'd4214;
		word[15'd5139] <= 32'd4215;
		word[15'd5140] <= 32'd4216;
		word[15'd5141] <= 32'd4217;
		word[15'd5142] <= 32'd4218;
		word[15'd5143] <= 32'd4219;
		word[15'd5144] <= 32'd4220;
		word[15'd5145] <= 32'd4221;
		word[15'd5146] <= 32'd4222;
		word[15'd5147] <= 32'd4223;
		word[15'd5148] <= 32'd4224;
		word[15'd5149] <= 32'd4225;
		word[15'd5150] <= 32'd4226;
		word[15'd5151] <= 32'd4227;
		word[15'd5152] <= 32'd4228;
		word[15'd5153] <= 32'd4229;
		word[15'd5154] <= 32'd4230;
		word[15'd5155] <= 32'd4231;
		word[15'd5156] <= 32'd4232;
		word[15'd5157] <= 32'd4233;
		word[15'd5158] <= 32'd4234;
		word[15'd5159] <= 32'd4235;
		word[15'd5160] <= 32'd4236;
		word[15'd5161] <= 32'd4237;
		word[15'd5162] <= 32'd4238;
		word[15'd5163] <= 32'd4239;
		word[15'd5164] <= 32'd4240;
		word[15'd5165] <= 32'd4241;
		word[15'd5166] <= 32'd4242;
		word[15'd5167] <= 32'd4243;
		word[15'd5168] <= 32'd4244;
		word[15'd5169] <= 32'd4245;
		word[15'd5170] <= 32'd4246;
		word[15'd5171] <= 32'd4247;
		word[15'd5172] <= 32'd4248;
		word[15'd5173] <= 32'd4249;
		word[15'd5174] <= 32'd4250;
		word[15'd5175] <= 32'd4251;
		word[15'd5176] <= 32'd4252;
		word[15'd5177] <= 32'd4253;
		word[15'd5178] <= 32'd4254;
		word[15'd5179] <= 32'd4255;
		word[15'd5180] <= 32'd4256;
		word[15'd5181] <= 32'd4257;
		word[15'd5182] <= 32'd4258;
		word[15'd5183] <= 32'd4259;
		word[15'd5184] <= 32'd4260;
		word[15'd5185] <= 32'd4261;
		word[15'd5186] <= 32'd4262;
		word[15'd5187] <= 32'd4263;
		word[15'd5188] <= 32'd4264;
		word[15'd5189] <= 32'd4265;
		word[15'd5190] <= 32'd4266;
		word[15'd5191] <= 32'd4267;
		word[15'd5192] <= 32'd4268;
		word[15'd5193] <= 32'd4269;
		word[15'd5194] <= 32'd4270;
		word[15'd5195] <= 32'd4271;
		word[15'd5196] <= 32'd4272;
		word[15'd5197] <= 32'd4273;
		word[15'd5198] <= 32'd4274;
		word[15'd5199] <= 32'd4275;
		word[15'd5200] <= 32'd4276;
		word[15'd5201] <= 32'd4277;
		word[15'd5202] <= 32'd4278;
		word[15'd5203] <= 32'd4279;
		word[15'd5204] <= 32'd4280;
		word[15'd5205] <= 32'd4281;
		word[15'd5206] <= 32'd4282;
		word[15'd5207] <= 32'd4283;
		word[15'd5208] <= 32'd4284;
		word[15'd5209] <= 32'd4285;
		word[15'd5210] <= 32'd4286;
		word[15'd5211] <= 32'd4287;
		word[15'd5212] <= 32'd4288;
		word[15'd5213] <= 32'd4289;
		word[15'd5214] <= 32'd4290;
		word[15'd5215] <= 32'd4291;
		word[15'd5216] <= 32'd4292;
		word[15'd5217] <= 32'd4293;
		word[15'd5218] <= 32'd4294;
		word[15'd5219] <= 32'd4295;
		word[15'd5220] <= 32'd4296;
		word[15'd5221] <= 32'd4297;
		word[15'd5222] <= 32'd4298;
		word[15'd5223] <= 32'd4299;
		word[15'd5224] <= 32'd4300;
		word[15'd5225] <= 32'd4301;
		word[15'd5226] <= 32'd4302;
		word[15'd5227] <= 32'd4303;
		word[15'd5228] <= 32'd4304;
		word[15'd5229] <= 32'd4305;
		word[15'd5230] <= 32'd4306;
		word[15'd5231] <= 32'd4307;
		word[15'd5232] <= 32'd4308;
		word[15'd5233] <= 32'd4309;
		word[15'd5234] <= 32'd4310;
		word[15'd5235] <= 32'd4311;
		word[15'd5236] <= 32'd4312;
		word[15'd5237] <= 32'd4313;
		word[15'd5238] <= 32'd4314;
		word[15'd5239] <= 32'd4315;
		word[15'd5240] <= 32'd4316;
		word[15'd5241] <= 32'd4317;
		word[15'd5242] <= 32'd4318;
		word[15'd5243] <= 32'd4319;
		word[15'd5244] <= 32'd4320;
		word[15'd5245] <= 32'd4321;
		word[15'd5246] <= 32'd4322;
		word[15'd5247] <= 32'd4323;
		word[15'd5248] <= 32'd4324;
		word[15'd5249] <= 32'd4325;
		word[15'd5250] <= 32'd4326;
		word[15'd5251] <= 32'd4327;
		word[15'd5252] <= 32'd4328;
		word[15'd5253] <= 32'd4329;
		word[15'd5254] <= 32'd4330;
		word[15'd5255] <= 32'd4331;
		word[15'd5256] <= 32'd4332;
		word[15'd5257] <= 32'd4333;
		word[15'd5258] <= 32'd4334;
		word[15'd5259] <= 32'd4335;
		word[15'd5260] <= 32'd4336;
		word[15'd5261] <= 32'd4337;
		word[15'd5262] <= 32'd4338;
		word[15'd5263] <= 32'd4339;
		word[15'd5264] <= 32'd4340;
		word[15'd5265] <= 32'd4341;
		word[15'd5266] <= 32'd4342;
		word[15'd5267] <= 32'd4343;
		word[15'd5268] <= 32'd4344;
		word[15'd5269] <= 32'd4345;
		word[15'd5270] <= 32'd4346;
		word[15'd5271] <= 32'd4347;
		word[15'd5272] <= 32'd4348;
		word[15'd5273] <= 32'd4349;
		word[15'd5274] <= 32'd4350;
		word[15'd5275] <= 32'd4351;
		word[15'd5276] <= 32'd4352;
		word[15'd5277] <= 32'd4353;
		word[15'd5278] <= 32'd4354;
		word[15'd5279] <= 32'd4355;
		word[15'd5280] <= 32'd4356;
		word[15'd5281] <= 32'd4357;
		word[15'd5282] <= 32'd4358;
		word[15'd5283] <= 32'd4359;
		word[15'd5284] <= 32'd4360;
		word[15'd5285] <= 32'd4361;
		word[15'd5286] <= 32'd4362;
		word[15'd5287] <= 32'd4363;
		word[15'd5288] <= 32'd4364;
		word[15'd5289] <= 32'd4365;
		word[15'd5290] <= 32'd4366;
		word[15'd5291] <= 32'd4367;
		word[15'd5292] <= 32'd4368;
		word[15'd5293] <= 32'd4369;
		word[15'd5294] <= 32'd4370;
		word[15'd5295] <= 32'd4371;
		word[15'd5296] <= 32'd4372;
		word[15'd5297] <= 32'd4373;
		word[15'd5298] <= 32'd4374;
		word[15'd5299] <= 32'd4375;
		word[15'd5300] <= 32'd4376;
		word[15'd5301] <= 32'd4377;
		word[15'd5302] <= 32'd4378;
		word[15'd5303] <= 32'd4379;
		word[15'd5304] <= 32'd4380;
		word[15'd5305] <= 32'd4381;
		word[15'd5306] <= 32'd4382;
		word[15'd5307] <= 32'd4383;
		word[15'd5308] <= 32'd4384;
		word[15'd5309] <= 32'd4385;
		word[15'd5310] <= 32'd4386;
		word[15'd5311] <= 32'd4387;
		word[15'd5312] <= 32'd4388;
		word[15'd5313] <= 32'd4389;
		word[15'd5314] <= 32'd4390;
		word[15'd5315] <= 32'd4391;
		word[15'd5316] <= 32'd4392;
		word[15'd5317] <= 32'd4393;
		word[15'd5318] <= 32'd4394;
		word[15'd5319] <= 32'd4395;
		word[15'd5320] <= 32'd4396;
		word[15'd5321] <= 32'd4397;
		word[15'd5322] <= 32'd4398;
		word[15'd5323] <= 32'd4399;
		word[15'd5324] <= 32'd4400;
		word[15'd5325] <= 32'd4401;
		word[15'd5326] <= 32'd4402;
		word[15'd5327] <= 32'd4403;
		word[15'd5328] <= 32'd4404;
		word[15'd5329] <= 32'd4405;
		word[15'd5330] <= 32'd4406;
		word[15'd5331] <= 32'd4407;
		word[15'd5332] <= 32'd4408;
		word[15'd5333] <= 32'd4409;
		word[15'd5334] <= 32'd4410;
		word[15'd5335] <= 32'd4411;
		word[15'd5336] <= 32'd4412;
		word[15'd5337] <= 32'd4413;
		word[15'd5338] <= 32'd4414;
		word[15'd5339] <= 32'd4415;
		word[15'd5340] <= 32'd4416;
		word[15'd5341] <= 32'd4417;
		word[15'd5342] <= 32'd4418;
		word[15'd5343] <= 32'd4419;
		word[15'd5344] <= 32'd4420;
		word[15'd5345] <= 32'd4421;
		word[15'd5346] <= 32'd4422;
		word[15'd5347] <= 32'd4423;
		word[15'd5348] <= 32'd4424;
		word[15'd5349] <= 32'd4425;
		word[15'd5350] <= 32'd4426;
		word[15'd5351] <= 32'd4427;
		word[15'd5352] <= 32'd4428;
		word[15'd5353] <= 32'd4429;
		word[15'd5354] <= 32'd4430;
		word[15'd5355] <= 32'd4431;
		word[15'd5356] <= 32'd4432;
		word[15'd5357] <= 32'd4433;
		word[15'd5358] <= 32'd4434;
		word[15'd5359] <= 32'd4435;
		word[15'd5360] <= 32'd4436;
		word[15'd5361] <= 32'd4437;
		word[15'd5362] <= 32'd4438;
		word[15'd5363] <= 32'd4439;
		word[15'd5364] <= 32'd4440;
		word[15'd5365] <= 32'd4441;
		word[15'd5366] <= 32'd4442;
		word[15'd5367] <= 32'd4443;
		word[15'd5368] <= 32'd4444;
		word[15'd5369] <= 32'd4445;
		word[15'd5370] <= 32'd4446;
		word[15'd5371] <= 32'd4447;
		word[15'd5372] <= 32'd4448;
		word[15'd5373] <= 32'd4449;
		word[15'd5374] <= 32'd4450;
		word[15'd5375] <= 32'd4451;
		word[15'd5376] <= 32'd4452;
		word[15'd5377] <= 32'd4453;
		word[15'd5378] <= 32'd4454;
		word[15'd5379] <= 32'd4455;
		word[15'd5380] <= 32'd4456;
		word[15'd5381] <= 32'd4457;
		word[15'd5382] <= 32'd4458;
		word[15'd5383] <= 32'd4459;
		word[15'd5384] <= 32'd4460;
		word[15'd5385] <= 32'd4461;
		word[15'd5386] <= 32'd4462;
		word[15'd5387] <= 32'd4463;
		word[15'd5388] <= 32'd4464;
		word[15'd5389] <= 32'd4465;
		word[15'd5390] <= 32'd4466;
		word[15'd5391] <= 32'd4467;
		word[15'd5392] <= 32'd4468;
		word[15'd5393] <= 32'd4469;
		word[15'd5394] <= 32'd4470;
		word[15'd5395] <= 32'd4471;
		word[15'd5396] <= 32'd4472;
		word[15'd5397] <= 32'd4473;
		word[15'd5398] <= 32'd4474;
		word[15'd5399] <= 32'd4475;
		word[15'd5400] <= 32'd4476;
		word[15'd5401] <= 32'd4477;
		word[15'd5402] <= 32'd4478;
		word[15'd5403] <= 32'd4479;
		word[15'd5404] <= 32'd4480;
		word[15'd5405] <= 32'd4481;
		word[15'd5406] <= 32'd4482;
		word[15'd5407] <= 32'd4483;
		word[15'd5408] <= 32'd4484;
		word[15'd5409] <= 32'd4485;
		word[15'd5410] <= 32'd4486;
		word[15'd5411] <= 32'd4487;
		word[15'd5412] <= 32'd4488;
		word[15'd5413] <= 32'd4489;
		word[15'd5414] <= 32'd4490;
		word[15'd5415] <= 32'd4491;
		word[15'd5416] <= 32'd4492;
		word[15'd5417] <= 32'd4493;
		word[15'd5418] <= 32'd4494;
		word[15'd5419] <= 32'd4495;
		word[15'd5420] <= 32'd4496;
		word[15'd5421] <= 32'd4497;
		word[15'd5422] <= 32'd4498;
		word[15'd5423] <= 32'd4499;
		word[15'd5424] <= 32'd4500;
		word[15'd5425] <= 32'd4501;
		word[15'd5426] <= 32'd4502;
		word[15'd5427] <= 32'd4503;
		word[15'd5428] <= 32'd4504;
		word[15'd5429] <= 32'd4505;
		word[15'd5430] <= 32'd4506;
		word[15'd5431] <= 32'd4507;
		word[15'd5432] <= 32'd4508;
		word[15'd5433] <= 32'd4509;
		word[15'd5434] <= 32'd4510;
		word[15'd5435] <= 32'd4511;
		word[15'd5436] <= 32'd4512;
		word[15'd5437] <= 32'd4513;
		word[15'd5438] <= 32'd4514;
		word[15'd5439] <= 32'd4515;
		word[15'd5440] <= 32'd4516;
		word[15'd5441] <= 32'd4517;
		word[15'd5442] <= 32'd4518;
		word[15'd5443] <= 32'd4519;
		word[15'd5444] <= 32'd4520;
		word[15'd5445] <= 32'd4521;
		word[15'd5446] <= 32'd4522;
		word[15'd5447] <= 32'd4523;
		word[15'd5448] <= 32'd4524;
		word[15'd5449] <= 32'd4525;
		word[15'd5450] <= 32'd4526;
		word[15'd5451] <= 32'd4527;
		word[15'd5452] <= 32'd4528;
		word[15'd5453] <= 32'd4529;
		word[15'd5454] <= 32'd4530;
		word[15'd5455] <= 32'd4531;
		word[15'd5456] <= 32'd4532;
		word[15'd5457] <= 32'd4533;
		word[15'd5458] <= 32'd4534;
		word[15'd5459] <= 32'd4535;
		word[15'd5460] <= 32'd4536;
		word[15'd5461] <= 32'd4537;
		word[15'd5462] <= 32'd4538;
		word[15'd5463] <= 32'd4539;
		word[15'd5464] <= 32'd4540;
		word[15'd5465] <= 32'd4541;
		word[15'd5466] <= 32'd4542;
		word[15'd5467] <= 32'd4543;
		word[15'd5468] <= 32'd4544;
		word[15'd5469] <= 32'd4545;
		word[15'd5470] <= 32'd4546;
		word[15'd5471] <= 32'd4547;
		word[15'd5472] <= 32'd4548;
		word[15'd5473] <= 32'd4549;
		word[15'd5474] <= 32'd4550;
		word[15'd5475] <= 32'd4551;
		word[15'd5476] <= 32'd4552;
		word[15'd5477] <= 32'd4553;
		word[15'd5478] <= 32'd4554;
		word[15'd5479] <= 32'd4555;
		word[15'd5480] <= 32'd4556;
		word[15'd5481] <= 32'd4557;
		word[15'd5482] <= 32'd4558;
		word[15'd5483] <= 32'd4559;
		word[15'd5484] <= 32'd4560;
		word[15'd5485] <= 32'd4561;
		word[15'd5486] <= 32'd4562;
		word[15'd5487] <= 32'd4563;
		word[15'd5488] <= 32'd4564;
		word[15'd5489] <= 32'd4565;
		word[15'd5490] <= 32'd4566;
		word[15'd5491] <= 32'd4567;
		word[15'd5492] <= 32'd4568;
		word[15'd5493] <= 32'd4569;
		word[15'd5494] <= 32'd4570;
		word[15'd5495] <= 32'd4571;
		word[15'd5496] <= 32'd4572;
		word[15'd5497] <= 32'd4573;
		word[15'd5498] <= 32'd4574;
		word[15'd5499] <= 32'd4575;
		word[15'd5500] <= 32'd4576;
		word[15'd5501] <= 32'd4577;
		word[15'd5502] <= 32'd4578;
		word[15'd5503] <= 32'd4579;
		word[15'd5504] <= 32'd4580;
		word[15'd5505] <= 32'd4581;
		word[15'd5506] <= 32'd4582;
		word[15'd5507] <= 32'd4583;
		word[15'd5508] <= 32'd4584;
		word[15'd5509] <= 32'd4585;
		word[15'd5510] <= 32'd4586;
		word[15'd5511] <= 32'd4587;
		word[15'd5512] <= 32'd4588;
		word[15'd5513] <= 32'd4589;
		word[15'd5514] <= 32'd4590;
		word[15'd5515] <= 32'd4591;
		word[15'd5516] <= 32'd4592;
		word[15'd5517] <= 32'd4593;
		word[15'd5518] <= 32'd4594;
		word[15'd5519] <= 32'd4595;
		word[15'd5520] <= 32'd4596;
		word[15'd5521] <= 32'd4597;
		word[15'd5522] <= 32'd4598;
		word[15'd5523] <= 32'd4599;
		word[15'd5524] <= 32'd4600;
		word[15'd5525] <= 32'd4601;
		word[15'd5526] <= 32'd4602;
		word[15'd5527] <= 32'd4603;
		word[15'd5528] <= 32'd4604;
		word[15'd5529] <= 32'd4605;
		word[15'd5530] <= 32'd4606;
		word[15'd5531] <= 32'd4607;
		word[15'd5532] <= 32'd4608;
		word[15'd5533] <= 32'd4609;
		word[15'd5534] <= 32'd4610;
		word[15'd5535] <= 32'd4611;
		word[15'd5536] <= 32'd4612;
		word[15'd5537] <= 32'd4613;
		word[15'd5538] <= 32'd4614;
		word[15'd5539] <= 32'd4615;
		word[15'd5540] <= 32'd4616;
		word[15'd5541] <= 32'd4617;
		word[15'd5542] <= 32'd4618;
		word[15'd5543] <= 32'd4619;
		word[15'd5544] <= 32'd4620;
		word[15'd5545] <= 32'd4621;
		word[15'd5546] <= 32'd4622;
		word[15'd5547] <= 32'd4623;
		word[15'd5548] <= 32'd4624;
		word[15'd5549] <= 32'd4625;
		word[15'd5550] <= 32'd4626;
		word[15'd5551] <= 32'd4627;
		word[15'd5552] <= 32'd4628;
		word[15'd5553] <= 32'd4629;
		word[15'd5554] <= 32'd4630;
		word[15'd5555] <= 32'd4631;
		word[15'd5556] <= 32'd4632;
		word[15'd5557] <= 32'd4633;
		word[15'd5558] <= 32'd4634;
		word[15'd5559] <= 32'd4635;
		word[15'd5560] <= 32'd4636;
		word[15'd5561] <= 32'd4637;
		word[15'd5562] <= 32'd4638;
		word[15'd5563] <= 32'd4639;
		word[15'd5564] <= 32'd4640;
		word[15'd5565] <= 32'd4641;
		word[15'd5566] <= 32'd4642;
		word[15'd5567] <= 32'd4643;
		word[15'd5568] <= 32'd4644;
		word[15'd5569] <= 32'd4645;
		word[15'd5570] <= 32'd4646;
		word[15'd5571] <= 32'd4647;
		word[15'd5572] <= 32'd4648;
		word[15'd5573] <= 32'd4649;
		word[15'd5574] <= 32'd4650;
		word[15'd5575] <= 32'd4651;
		word[15'd5576] <= 32'd4652;
		word[15'd5577] <= 32'd4653;
		word[15'd5578] <= 32'd4654;
		word[15'd5579] <= 32'd4655;
		word[15'd5580] <= 32'd4656;
		word[15'd5581] <= 32'd4657;
		word[15'd5582] <= 32'd4658;
		word[15'd5583] <= 32'd4659;
		word[15'd5584] <= 32'd4660;
		word[15'd5585] <= 32'd4661;
		word[15'd5586] <= 32'd4662;
		word[15'd5587] <= 32'd4663;
		word[15'd5588] <= 32'd4664;
		word[15'd5589] <= 32'd4665;
		word[15'd5590] <= 32'd4666;
		word[15'd5591] <= 32'd4667;
		word[15'd5592] <= 32'd4668;
		word[15'd5593] <= 32'd4669;
		word[15'd5594] <= 32'd4670;
		word[15'd5595] <= 32'd4671;
		word[15'd5596] <= 32'd4672;
		word[15'd5597] <= 32'd4673;
		word[15'd5598] <= 32'd4674;
		word[15'd5599] <= 32'd4675;
		word[15'd5600] <= 32'd4676;
		word[15'd5601] <= 32'd4677;
		word[15'd5602] <= 32'd4678;
		word[15'd5603] <= 32'd4679;
		word[15'd5604] <= 32'd4680;
		word[15'd5605] <= 32'd4681;
		word[15'd5606] <= 32'd4682;
		word[15'd5607] <= 32'd4683;
		word[15'd5608] <= 32'd4684;
		word[15'd5609] <= 32'd4685;
		word[15'd5610] <= 32'd4686;
		word[15'd5611] <= 32'd4687;
		word[15'd5612] <= 32'd4688;
		word[15'd5613] <= 32'd4689;
		word[15'd5614] <= 32'd4690;
		word[15'd5615] <= 32'd4691;
		word[15'd5616] <= 32'd4692;
		word[15'd5617] <= 32'd4693;
		word[15'd5618] <= 32'd4694;
		word[15'd5619] <= 32'd4695;
		word[15'd5620] <= 32'd4696;
		word[15'd5621] <= 32'd4697;
		word[15'd5622] <= 32'd4698;
		word[15'd5623] <= 32'd4699;
		word[15'd5624] <= 32'd4700;
		word[15'd5625] <= 32'd4701;
		word[15'd5626] <= 32'd4702;
		word[15'd5627] <= 32'd4703;
		word[15'd5628] <= 32'd4704;
		word[15'd5629] <= 32'd4705;
		word[15'd5630] <= 32'd4706;
		word[15'd5631] <= 32'd4707;
		word[15'd5632] <= 32'd4708;
		word[15'd5633] <= 32'd4709;
		word[15'd5634] <= 32'd4710;
		word[15'd5635] <= 32'd4711;
		word[15'd5636] <= 32'd4712;
		word[15'd5637] <= 32'd4713;
		word[15'd5638] <= 32'd4714;
		word[15'd5639] <= 32'd4715;
		word[15'd5640] <= 32'd4716;
		word[15'd5641] <= 32'd4717;
		word[15'd5642] <= 32'd4718;
		word[15'd5643] <= 32'd4719;
		word[15'd5644] <= 32'd4720;
		word[15'd5645] <= 32'd4721;
		word[15'd5646] <= 32'd4722;
		word[15'd5647] <= 32'd4723;
		word[15'd5648] <= 32'd4724;
		word[15'd5649] <= 32'd4725;
		word[15'd5650] <= 32'd4726;
		word[15'd5651] <= 32'd4727;
		word[15'd5652] <= 32'd4728;
		word[15'd5653] <= 32'd4729;
		word[15'd5654] <= 32'd4730;
		word[15'd5655] <= 32'd4731;
		word[15'd5656] <= 32'd4732;
		word[15'd5657] <= 32'd4733;
		word[15'd5658] <= 32'd4734;
		word[15'd5659] <= 32'd4735;
		word[15'd5660] <= 32'd4736;
		word[15'd5661] <= 32'd4737;
		word[15'd5662] <= 32'd4738;
		word[15'd5663] <= 32'd4739;
		word[15'd5664] <= 32'd4740;
		word[15'd5665] <= 32'd4741;
		word[15'd5666] <= 32'd4742;
		word[15'd5667] <= 32'd4743;
		word[15'd5668] <= 32'd4744;
		word[15'd5669] <= 32'd4745;
		word[15'd5670] <= 32'd4746;
		word[15'd5671] <= 32'd4747;
		word[15'd5672] <= 32'd4748;
		word[15'd5673] <= 32'd4749;
		word[15'd5674] <= 32'd4750;
		word[15'd5675] <= 32'd4751;
		word[15'd5676] <= 32'd4752;
		word[15'd5677] <= 32'd4753;
		word[15'd5678] <= 32'd4754;
		word[15'd5679] <= 32'd4755;
		word[15'd5680] <= 32'd4756;
		word[15'd5681] <= 32'd4757;
		word[15'd5682] <= 32'd4758;
		word[15'd5683] <= 32'd4759;
		word[15'd5684] <= 32'd4760;
		word[15'd5685] <= 32'd4761;
		word[15'd5686] <= 32'd4762;
		word[15'd5687] <= 32'd4763;
		word[15'd5688] <= 32'd4764;
		word[15'd5689] <= 32'd4765;
		word[15'd5690] <= 32'd4766;
		word[15'd5691] <= 32'd4767;
		word[15'd5692] <= 32'd4768;
		word[15'd5693] <= 32'd4769;
		word[15'd5694] <= 32'd4770;
		word[15'd5695] <= 32'd4771;
		word[15'd5696] <= 32'd4772;
		word[15'd5697] <= 32'd4773;
		word[15'd5698] <= 32'd4774;
		word[15'd5699] <= 32'd4775;
		word[15'd5700] <= 32'd4776;
		word[15'd5701] <= 32'd4777;
		word[15'd5702] <= 32'd4778;
		word[15'd5703] <= 32'd4779;
		word[15'd5704] <= 32'd4780;
		word[15'd5705] <= 32'd4781;
		word[15'd5706] <= 32'd4782;
		word[15'd5707] <= 32'd4783;
		word[15'd5708] <= 32'd4784;
		word[15'd5709] <= 32'd4785;
		word[15'd5710] <= 32'd4786;
		word[15'd5711] <= 32'd4787;
		word[15'd5712] <= 32'd4788;
		word[15'd5713] <= 32'd4789;
		word[15'd5714] <= 32'd4790;
		word[15'd5715] <= 32'd4791;
		word[15'd5716] <= 32'd4792;
		word[15'd5717] <= 32'd4793;
		word[15'd5718] <= 32'd4794;
		word[15'd5719] <= 32'd4795;
		word[15'd5720] <= 32'd4796;
		word[15'd5721] <= 32'd4797;
		word[15'd5722] <= 32'd4798;
		word[15'd5723] <= 32'd4799;
		word[15'd5724] <= 32'd4800;
		word[15'd5725] <= 32'd4801;
		word[15'd5726] <= 32'd4802;
		word[15'd5727] <= 32'd4803;
		word[15'd5728] <= 32'd4804;
		word[15'd5729] <= 32'd4805;
		word[15'd5730] <= 32'd4806;
		word[15'd5731] <= 32'd4807;
		word[15'd5732] <= 32'd4808;
		word[15'd5733] <= 32'd4809;
		word[15'd5734] <= 32'd4810;
		word[15'd5735] <= 32'd4811;
		word[15'd5736] <= 32'd4812;
		word[15'd5737] <= 32'd4813;
		word[15'd5738] <= 32'd4814;
		word[15'd5739] <= 32'd4815;
		word[15'd5740] <= 32'd4816;
		word[15'd5741] <= 32'd4817;
		word[15'd5742] <= 32'd4818;
		word[15'd5743] <= 32'd4819;
		word[15'd5744] <= 32'd4820;
		word[15'd5745] <= 32'd4821;
		word[15'd5746] <= 32'd4822;
		word[15'd5747] <= 32'd4823;
		word[15'd5748] <= 32'd4824;
		word[15'd5749] <= 32'd4825;
		word[15'd5750] <= 32'd4826;
		word[15'd5751] <= 32'd4827;
		word[15'd5752] <= 32'd4828;
		word[15'd5753] <= 32'd4829;
		word[15'd5754] <= 32'd4830;
		word[15'd5755] <= 32'd4831;
		word[15'd5756] <= 32'd4832;
		word[15'd5757] <= 32'd4833;
		word[15'd5758] <= 32'd4834;
		word[15'd5759] <= 32'd4835;
		word[15'd5760] <= 32'd4836;
		word[15'd5761] <= 32'd4837;
		word[15'd5762] <= 32'd4838;
		word[15'd5763] <= 32'd4839;
		word[15'd5764] <= 32'd4840;
		word[15'd5765] <= 32'd4841;
		word[15'd5766] <= 32'd4842;
		word[15'd5767] <= 32'd4843;
		word[15'd5768] <= 32'd4844;
		word[15'd5769] <= 32'd4845;
		word[15'd5770] <= 32'd4846;
		word[15'd5771] <= 32'd4847;
		word[15'd5772] <= 32'd4848;
		word[15'd5773] <= 32'd4849;
		word[15'd5774] <= 32'd4850;
		word[15'd5775] <= 32'd4851;
		word[15'd5776] <= 32'd4852;
		word[15'd5777] <= 32'd4853;
		word[15'd5778] <= 32'd4854;
		word[15'd5779] <= 32'd4855;
		word[15'd5780] <= 32'd4856;
		word[15'd5781] <= 32'd4857;
		word[15'd5782] <= 32'd4858;
		word[15'd5783] <= 32'd4859;
		word[15'd5784] <= 32'd4860;
		word[15'd5785] <= 32'd4861;
		word[15'd5786] <= 32'd4862;
		word[15'd5787] <= 32'd4863;
		word[15'd5788] <= 32'd4864;
		word[15'd5789] <= 32'd4865;
		word[15'd5790] <= 32'd4866;
		word[15'd5791] <= 32'd4867;
		word[15'd5792] <= 32'd4868;
		word[15'd5793] <= 32'd4869;
		word[15'd5794] <= 32'd4870;
		word[15'd5795] <= 32'd4871;
		word[15'd5796] <= 32'd4872;
		word[15'd5797] <= 32'd4873;
		word[15'd5798] <= 32'd4874;
		word[15'd5799] <= 32'd4875;
		word[15'd5800] <= 32'd4876;
		word[15'd5801] <= 32'd4877;
		word[15'd5802] <= 32'd4878;
		word[15'd5803] <= 32'd4879;
		word[15'd5804] <= 32'd4880;
		word[15'd5805] <= 32'd4881;
		word[15'd5806] <= 32'd4882;
		word[15'd5807] <= 32'd4883;
		word[15'd5808] <= 32'd4884;
		word[15'd5809] <= 32'd4885;
		word[15'd5810] <= 32'd4886;
		word[15'd5811] <= 32'd4887;
		word[15'd5812] <= 32'd4888;
		word[15'd5813] <= 32'd4889;
		word[15'd5814] <= 32'd4890;
		word[15'd5815] <= 32'd4891;
		word[15'd5816] <= 32'd4892;
		word[15'd5817] <= 32'd4893;
		word[15'd5818] <= 32'd4894;
		word[15'd5819] <= 32'd4895;
		word[15'd5820] <= 32'd4896;
		word[15'd5821] <= 32'd4897;
		word[15'd5822] <= 32'd4898;
		word[15'd5823] <= 32'd4899;
		word[15'd5824] <= 32'd4900;
		word[15'd5825] <= 32'd4901;
		word[15'd5826] <= 32'd4902;
		word[15'd5827] <= 32'd4903;
		word[15'd5828] <= 32'd4904;
		word[15'd5829] <= 32'd4905;
		word[15'd5830] <= 32'd4906;
		word[15'd5831] <= 32'd4907;
		word[15'd5832] <= 32'd4908;
		word[15'd5833] <= 32'd4909;
		word[15'd5834] <= 32'd4910;
		word[15'd5835] <= 32'd4911;
		word[15'd5836] <= 32'd4912;
		word[15'd5837] <= 32'd4913;
		word[15'd5838] <= 32'd4914;
		word[15'd5839] <= 32'd4915;
		word[15'd5840] <= 32'd4916;
		word[15'd5841] <= 32'd4917;
		word[15'd5842] <= 32'd4918;
		word[15'd5843] <= 32'd4919;
		word[15'd5844] <= 32'd4920;
		word[15'd5845] <= 32'd4921;
		word[15'd5846] <= 32'd4922;
		word[15'd5847] <= 32'd4923;
		word[15'd5848] <= 32'd4924;
		word[15'd5849] <= 32'd4925;
		word[15'd5850] <= 32'd4926;
		word[15'd5851] <= 32'd4927;
		word[15'd5852] <= 32'd4928;
		word[15'd5853] <= 32'd4929;
		word[15'd5854] <= 32'd4930;
		word[15'd5855] <= 32'd4931;
		word[15'd5856] <= 32'd4932;
		word[15'd5857] <= 32'd4933;
		word[15'd5858] <= 32'd4934;
		word[15'd5859] <= 32'd4935;
		word[15'd5860] <= 32'd4936;
		word[15'd5861] <= 32'd4937;
		word[15'd5862] <= 32'd4938;
		word[15'd5863] <= 32'd4939;
		word[15'd5864] <= 32'd4940;
		word[15'd5865] <= 32'd4941;
		word[15'd5866] <= 32'd4942;
		word[15'd5867] <= 32'd4943;
		word[15'd5868] <= 32'd4944;
		word[15'd5869] <= 32'd4945;
		word[15'd5870] <= 32'd4946;
		word[15'd5871] <= 32'd4947;
		word[15'd5872] <= 32'd4948;
		word[15'd5873] <= 32'd4949;
		word[15'd5874] <= 32'd4950;
		word[15'd5875] <= 32'd4951;
		word[15'd5876] <= 32'd4952;
		word[15'd5877] <= 32'd4953;
		word[15'd5878] <= 32'd4954;
		word[15'd5879] <= 32'd4955;
		word[15'd5880] <= 32'd4956;
		word[15'd5881] <= 32'd4957;
		word[15'd5882] <= 32'd4958;
		word[15'd5883] <= 32'd4959;
		word[15'd5884] <= 32'd4960;
		word[15'd5885] <= 32'd4961;
		word[15'd5886] <= 32'd4962;
		word[15'd5887] <= 32'd4963;
		word[15'd5888] <= 32'd4964;
		word[15'd5889] <= 32'd4965;
		word[15'd5890] <= 32'd4966;
		word[15'd5891] <= 32'd4967;
		word[15'd5892] <= 32'd4968;
		word[15'd5893] <= 32'd4969;
		word[15'd5894] <= 32'd4970;
		word[15'd5895] <= 32'd4971;
		word[15'd5896] <= 32'd4972;
		word[15'd5897] <= 32'd4973;
		word[15'd5898] <= 32'd4974;
		word[15'd5899] <= 32'd4975;
		word[15'd5900] <= 32'd4976;
		word[15'd5901] <= 32'd4977;
		word[15'd5902] <= 32'd4978;
		word[15'd5903] <= 32'd4979;
		word[15'd5904] <= 32'd4980;
		word[15'd5905] <= 32'd4981;
		word[15'd5906] <= 32'd4982;
		word[15'd5907] <= 32'd4983;
		word[15'd5908] <= 32'd4984;
		word[15'd5909] <= 32'd4985;
		word[15'd5910] <= 32'd4986;
		word[15'd5911] <= 32'd4987;
		word[15'd5912] <= 32'd4988;
		word[15'd5913] <= 32'd4989;
		word[15'd5914] <= 32'd4990;
		word[15'd5915] <= 32'd4991;
		word[15'd5916] <= 32'd4992;
		word[15'd5917] <= 32'd4993;
		word[15'd5918] <= 32'd4994;
		word[15'd5919] <= 32'd4995;
		word[15'd5920] <= 32'd4996;
		word[15'd5921] <= 32'd4997;
		word[15'd5922] <= 32'd4998;
		word[15'd5923] <= 32'd4999;
		word[15'd5924] <= 32'd5000;
		word[15'd5925] <= 32'd5001;
		word[15'd5926] <= 32'd5002;
		word[15'd5927] <= 32'd5003;
		word[15'd5928] <= 32'd5004;
		word[15'd5929] <= 32'd5005;
		word[15'd5930] <= 32'd5006;
		word[15'd5931] <= 32'd5007;
		word[15'd5932] <= 32'd5008;
		word[15'd5933] <= 32'd5009;
		word[15'd5934] <= 32'd5010;
		word[15'd5935] <= 32'd5011;
		word[15'd5936] <= 32'd5012;
		word[15'd5937] <= 32'd5013;
		word[15'd5938] <= 32'd5014;
		word[15'd5939] <= 32'd5015;
		word[15'd5940] <= 32'd5016;
		word[15'd5941] <= 32'd5017;
		word[15'd5942] <= 32'd5018;
		word[15'd5943] <= 32'd5019;
		word[15'd5944] <= 32'd5020;
		word[15'd5945] <= 32'd5021;
		word[15'd5946] <= 32'd5022;
		word[15'd5947] <= 32'd5023;
		word[15'd5948] <= 32'd5024;
		word[15'd5949] <= 32'd5025;
		word[15'd5950] <= 32'd5026;
		word[15'd5951] <= 32'd5027;
		word[15'd5952] <= 32'd5028;
		word[15'd5953] <= 32'd5029;
		word[15'd5954] <= 32'd5030;
		word[15'd5955] <= 32'd5031;
		word[15'd5956] <= 32'd5032;
		word[15'd5957] <= 32'd5033;
		word[15'd5958] <= 32'd5034;
		word[15'd5959] <= 32'd5035;
		word[15'd5960] <= 32'd5036;
		word[15'd5961] <= 32'd5037;
		word[15'd5962] <= 32'd5038;
		word[15'd5963] <= 32'd5039;
		word[15'd5964] <= 32'd5040;
		word[15'd5965] <= 32'd5041;
		word[15'd5966] <= 32'd5042;
		word[15'd5967] <= 32'd5043;
		word[15'd5968] <= 32'd5044;
		word[15'd5969] <= 32'd5045;
		word[15'd5970] <= 32'd5046;
		word[15'd5971] <= 32'd5047;
		word[15'd5972] <= 32'd5048;
		word[15'd5973] <= 32'd5049;
		word[15'd5974] <= 32'd5050;
		word[15'd5975] <= 32'd5051;
		word[15'd5976] <= 32'd5052;
		word[15'd5977] <= 32'd5053;
		word[15'd5978] <= 32'd5054;
		word[15'd5979] <= 32'd5055;
		word[15'd5980] <= 32'd5056;
		word[15'd5981] <= 32'd5057;
		word[15'd5982] <= 32'd5058;
		word[15'd5983] <= 32'd5059;
		word[15'd5984] <= 32'd5060;
		word[15'd5985] <= 32'd5061;
		word[15'd5986] <= 32'd5062;
		word[15'd5987] <= 32'd5063;
		word[15'd5988] <= 32'd5064;
		word[15'd5989] <= 32'd5065;
		word[15'd5990] <= 32'd5066;
		word[15'd5991] <= 32'd5067;
		word[15'd5992] <= 32'd5068;
		word[15'd5993] <= 32'd5069;
		word[15'd5994] <= 32'd5070;
		word[15'd5995] <= 32'd5071;
		word[15'd5996] <= 32'd5072;
		word[15'd5997] <= 32'd5073;
		word[15'd5998] <= 32'd5074;
		word[15'd5999] <= 32'd5075;
		word[15'd6000] <= 32'd5076;
		word[15'd6001] <= 32'd5077;
		word[15'd6002] <= 32'd5078;
		word[15'd6003] <= 32'd5079;
		word[15'd6004] <= 32'd5080;
		word[15'd6005] <= 32'd5081;
		word[15'd6006] <= 32'd5082;
		word[15'd6007] <= 32'd5083;
		word[15'd6008] <= 32'd5084;
		word[15'd6009] <= 32'd5085;
		word[15'd6010] <= 32'd5086;
		word[15'd6011] <= 32'd5087;
		word[15'd6012] <= 32'd5088;
		word[15'd6013] <= 32'd5089;
		word[15'd6014] <= 32'd5090;
		word[15'd6015] <= 32'd5091;
		word[15'd6016] <= 32'd5092;
		word[15'd6017] <= 32'd5093;
		word[15'd6018] <= 32'd5094;
		word[15'd6019] <= 32'd5095;
		word[15'd6020] <= 32'd5096;
		word[15'd6021] <= 32'd5097;
		word[15'd6022] <= 32'd5098;
		word[15'd6023] <= 32'd5099;
		word[15'd6024] <= 32'd5100;
		word[15'd6025] <= 32'd5101;
		word[15'd6026] <= 32'd5102;
		word[15'd6027] <= 32'd5103;
		word[15'd6028] <= 32'd5104;
		word[15'd6029] <= 32'd5105;
		word[15'd6030] <= 32'd5106;
		word[15'd6031] <= 32'd5107;
		word[15'd6032] <= 32'd5108;
		word[15'd6033] <= 32'd5109;
		word[15'd6034] <= 32'd5110;
		word[15'd6035] <= 32'd5111;
		word[15'd6036] <= 32'd5112;
		word[15'd6037] <= 32'd5113;
		word[15'd6038] <= 32'd5114;
		word[15'd6039] <= 32'd5115;
		word[15'd6040] <= 32'd5116;
		word[15'd6041] <= 32'd5117;
		word[15'd6042] <= 32'd5118;
		word[15'd6043] <= 32'd5119;
		word[15'd6044] <= 32'd5120;
		word[15'd6045] <= 32'd5121;
		word[15'd6046] <= 32'd5122;
		word[15'd6047] <= 32'd5123;
		word[15'd6048] <= 32'd5124;
		word[15'd6049] <= 32'd5125;
		word[15'd6050] <= 32'd5126;
		word[15'd6051] <= 32'd5127;
		word[15'd6052] <= 32'd5128;
		word[15'd6053] <= 32'd5129;
		word[15'd6054] <= 32'd5130;
		word[15'd6055] <= 32'd5131;
		word[15'd6056] <= 32'd5132;
		word[15'd6057] <= 32'd5133;
		word[15'd6058] <= 32'd5134;
		word[15'd6059] <= 32'd5135;
		word[15'd6060] <= 32'd5136;
		word[15'd6061] <= 32'd5137;
		word[15'd6062] <= 32'd5138;
		word[15'd6063] <= 32'd5139;
		word[15'd6064] <= 32'd5140;
		word[15'd6065] <= 32'd5141;
		word[15'd6066] <= 32'd5142;
		word[15'd6067] <= 32'd5143;
		word[15'd6068] <= 32'd5144;
		word[15'd6069] <= 32'd5145;
		word[15'd6070] <= 32'd5146;
		word[15'd6071] <= 32'd5147;
		word[15'd6072] <= 32'd5148;
		word[15'd6073] <= 32'd5149;
		word[15'd6074] <= 32'd5150;
		word[15'd6075] <= 32'd5151;
		word[15'd6076] <= 32'd5152;
		word[15'd6077] <= 32'd5153;
		word[15'd6078] <= 32'd5154;
		word[15'd6079] <= 32'd5155;
		word[15'd6080] <= 32'd5156;
		word[15'd6081] <= 32'd5157;
		word[15'd6082] <= 32'd5158;
		word[15'd6083] <= 32'd5159;
		word[15'd6084] <= 32'd5160;
		word[15'd6085] <= 32'd5161;
		word[15'd6086] <= 32'd5162;
		word[15'd6087] <= 32'd5163;
		word[15'd6088] <= 32'd5164;
		word[15'd6089] <= 32'd5165;
		word[15'd6090] <= 32'd5166;
		word[15'd6091] <= 32'd5167;
		word[15'd6092] <= 32'd5168;
		word[15'd6093] <= 32'd5169;
		word[15'd6094] <= 32'd5170;
		word[15'd6095] <= 32'd5171;
		word[15'd6096] <= 32'd5172;
		word[15'd6097] <= 32'd5173;
		word[15'd6098] <= 32'd5174;
		word[15'd6099] <= 32'd5175;
		word[15'd6100] <= 32'd5176;
		word[15'd6101] <= 32'd5177;
		word[15'd6102] <= 32'd5178;
		word[15'd6103] <= 32'd5179;
		word[15'd6104] <= 32'd5180;
		word[15'd6105] <= 32'd5181;
		word[15'd6106] <= 32'd5182;
		word[15'd6107] <= 32'd5183;
		word[15'd6108] <= 32'd5184;
		word[15'd6109] <= 32'd5185;
		word[15'd6110] <= 32'd5186;
		word[15'd6111] <= 32'd5187;
		word[15'd6112] <= 32'd5188;
		word[15'd6113] <= 32'd5189;
		word[15'd6114] <= 32'd5190;
		word[15'd6115] <= 32'd5191;
		word[15'd6116] <= 32'd5192;
		word[15'd6117] <= 32'd5193;
		word[15'd6118] <= 32'd5194;
		word[15'd6119] <= 32'd5195;
		word[15'd6120] <= 32'd5196;
		word[15'd6121] <= 32'd5197;
		word[15'd6122] <= 32'd5198;
		word[15'd6123] <= 32'd5199;
		word[15'd6124] <= 32'd5200;
		word[15'd6125] <= 32'd5201;
		word[15'd6126] <= 32'd5202;
		word[15'd6127] <= 32'd5203;
		word[15'd6128] <= 32'd5204;
		word[15'd6129] <= 32'd5205;
		word[15'd6130] <= 32'd5206;
		word[15'd6131] <= 32'd5207;
		word[15'd6132] <= 32'd5208;
		word[15'd6133] <= 32'd5209;
		word[15'd6134] <= 32'd5210;
		word[15'd6135] <= 32'd5211;
		word[15'd6136] <= 32'd5212;
		word[15'd6137] <= 32'd5213;
		word[15'd6138] <= 32'd5214;
		word[15'd6139] <= 32'd5215;
		word[15'd6140] <= 32'd5216;
		word[15'd6141] <= 32'd5217;
		word[15'd6142] <= 32'd5218;
		word[15'd6143] <= 32'd5219;
		word[15'd6144] <= 32'd5220;
		word[15'd6145] <= 32'd5221;
		word[15'd6146] <= 32'd5222;
		word[15'd6147] <= 32'd5223;
		word[15'd6148] <= 32'd5224;
		word[15'd6149] <= 32'd5225;
		word[15'd6150] <= 32'd5226;
		word[15'd6151] <= 32'd5227;
		word[15'd6152] <= 32'd5228;
		word[15'd6153] <= 32'd5229;
		word[15'd6154] <= 32'd5230;
		word[15'd6155] <= 32'd5231;
		word[15'd6156] <= 32'd5232;
		word[15'd6157] <= 32'd5233;
		word[15'd6158] <= 32'd5234;
		word[15'd6159] <= 32'd5235;
		word[15'd6160] <= 32'd5236;
		word[15'd6161] <= 32'd5237;
		word[15'd6162] <= 32'd5238;
		word[15'd6163] <= 32'd5239;
		word[15'd6164] <= 32'd5240;
		word[15'd6165] <= 32'd5241;
		word[15'd6166] <= 32'd5242;
		word[15'd6167] <= 32'd5243;
		word[15'd6168] <= 32'd5244;
		word[15'd6169] <= 32'd5245;
		word[15'd6170] <= 32'd5246;
		word[15'd6171] <= 32'd5247;
		word[15'd6172] <= 32'd5248;
		word[15'd6173] <= 32'd5249;
		word[15'd6174] <= 32'd5250;
		word[15'd6175] <= 32'd5251;
		word[15'd6176] <= 32'd5252;
		word[15'd6177] <= 32'd5253;
		word[15'd6178] <= 32'd5254;
		word[15'd6179] <= 32'd5255;
		word[15'd6180] <= 32'd5256;
		word[15'd6181] <= 32'd5257;
		word[15'd6182] <= 32'd5258;
		word[15'd6183] <= 32'd5259;
		word[15'd6184] <= 32'd5260;
		word[15'd6185] <= 32'd5261;
		word[15'd6186] <= 32'd5262;
		word[15'd6187] <= 32'd5263;
		word[15'd6188] <= 32'd5264;
		word[15'd6189] <= 32'd5265;
		word[15'd6190] <= 32'd5266;
		word[15'd6191] <= 32'd5267;
		word[15'd6192] <= 32'd5268;
		word[15'd6193] <= 32'd5269;
		word[15'd6194] <= 32'd5270;
		word[15'd6195] <= 32'd5271;
		word[15'd6196] <= 32'd5272;
		word[15'd6197] <= 32'd5273;
		word[15'd6198] <= 32'd5274;
		word[15'd6199] <= 32'd5275;
		word[15'd6200] <= 32'd5276;
		word[15'd6201] <= 32'd5277;
		word[15'd6202] <= 32'd5278;
		word[15'd6203] <= 32'd5279;
		word[15'd6204] <= 32'd5280;
		word[15'd6205] <= 32'd5281;
		word[15'd6206] <= 32'd5282;
		word[15'd6207] <= 32'd5283;
		word[15'd6208] <= 32'd5284;
		word[15'd6209] <= 32'd5285;
		word[15'd6210] <= 32'd5286;
		word[15'd6211] <= 32'd5287;
		word[15'd6212] <= 32'd5288;
		word[15'd6213] <= 32'd5289;
		word[15'd6214] <= 32'd5290;
		word[15'd6215] <= 32'd5291;
		word[15'd6216] <= 32'd5292;
		word[15'd6217] <= 32'd5293;
		word[15'd6218] <= 32'd5294;
		word[15'd6219] <= 32'd5295;
		word[15'd6220] <= 32'd5296;
		word[15'd6221] <= 32'd5297;
		word[15'd6222] <= 32'd5298;
		word[15'd6223] <= 32'd5299;
		word[15'd6224] <= 32'd5300;
		word[15'd6225] <= 32'd5301;
		word[15'd6226] <= 32'd5302;
		word[15'd6227] <= 32'd5303;
		word[15'd6228] <= 32'd5304;
		word[15'd6229] <= 32'd5305;
		word[15'd6230] <= 32'd5306;
		word[15'd6231] <= 32'd5307;
		word[15'd6232] <= 32'd5308;
		word[15'd6233] <= 32'd5309;
		word[15'd6234] <= 32'd5310;
		word[15'd6235] <= 32'd5311;
		word[15'd6236] <= 32'd5312;
		word[15'd6237] <= 32'd5313;
		word[15'd6238] <= 32'd5314;
		word[15'd6239] <= 32'd5315;
		word[15'd6240] <= 32'd5316;
		word[15'd6241] <= 32'd5317;
		word[15'd6242] <= 32'd5318;
		word[15'd6243] <= 32'd5319;
		word[15'd6244] <= 32'd5320;
		word[15'd6245] <= 32'd5321;
		word[15'd6246] <= 32'd5322;
		word[15'd6247] <= 32'd5323;
		word[15'd6248] <= 32'd5324;
		word[15'd6249] <= 32'd5325;
		word[15'd6250] <= 32'd5326;
		word[15'd6251] <= 32'd5327;
		word[15'd6252] <= 32'd5328;
		word[15'd6253] <= 32'd5329;
		word[15'd6254] <= 32'd5330;
		word[15'd6255] <= 32'd5331;
		word[15'd6256] <= 32'd5332;
		word[15'd6257] <= 32'd5333;
		word[15'd6258] <= 32'd5334;
		word[15'd6259] <= 32'd5335;
		word[15'd6260] <= 32'd5336;
		word[15'd6261] <= 32'd5337;
		word[15'd6262] <= 32'd5338;
		word[15'd6263] <= 32'd5339;
		word[15'd6264] <= 32'd5340;
		word[15'd6265] <= 32'd5341;
		word[15'd6266] <= 32'd5342;
		word[15'd6267] <= 32'd5343;
		word[15'd6268] <= 32'd5344;
		word[15'd6269] <= 32'd5345;
		word[15'd6270] <= 32'd5346;
		word[15'd6271] <= 32'd5347;
		word[15'd6272] <= 32'd5348;
		word[15'd6273] <= 32'd5349;
		word[15'd6274] <= 32'd5350;
		word[15'd6275] <= 32'd5351;
		word[15'd6276] <= 32'd5352;
		word[15'd6277] <= 32'd5353;
		word[15'd6278] <= 32'd5354;
		word[15'd6279] <= 32'd5355;
		word[15'd6280] <= 32'd5356;
		word[15'd6281] <= 32'd5357;
		word[15'd6282] <= 32'd5358;
		word[15'd6283] <= 32'd5359;
		word[15'd6284] <= 32'd5360;
		word[15'd6285] <= 32'd5361;
		word[15'd6286] <= 32'd5362;
		word[15'd6287] <= 32'd5363;
		word[15'd6288] <= 32'd5364;
		word[15'd6289] <= 32'd5365;
		word[15'd6290] <= 32'd5366;
		word[15'd6291] <= 32'd5367;
		word[15'd6292] <= 32'd5368;
		word[15'd6293] <= 32'd5369;
		word[15'd6294] <= 32'd5370;
		word[15'd6295] <= 32'd5371;
		word[15'd6296] <= 32'd5372;
		word[15'd6297] <= 32'd5373;
		word[15'd6298] <= 32'd5374;
		word[15'd6299] <= 32'd5375;
		word[15'd6300] <= 32'd5376;
		word[15'd6301] <= 32'd5377;
		word[15'd6302] <= 32'd5378;
		word[15'd6303] <= 32'd5379;
		word[15'd6304] <= 32'd5380;
		word[15'd6305] <= 32'd5381;
		word[15'd6306] <= 32'd5382;
		word[15'd6307] <= 32'd5383;
		word[15'd6308] <= 32'd5384;
		word[15'd6309] <= 32'd5385;
		word[15'd6310] <= 32'd5386;
		word[15'd6311] <= 32'd5387;
		word[15'd6312] <= 32'd5388;
		word[15'd6313] <= 32'd5389;
		word[15'd6314] <= 32'd5390;
		word[15'd6315] <= 32'd5391;
		word[15'd6316] <= 32'd5392;
		word[15'd6317] <= 32'd5393;
		word[15'd6318] <= 32'd5394;
		word[15'd6319] <= 32'd5395;
		word[15'd6320] <= 32'd5396;
		word[15'd6321] <= 32'd5397;
		word[15'd6322] <= 32'd5398;
		word[15'd6323] <= 32'd5399;
		word[15'd6324] <= 32'd5400;
		word[15'd6325] <= 32'd5401;
		word[15'd6326] <= 32'd5402;
		word[15'd6327] <= 32'd5403;
		word[15'd6328] <= 32'd5404;
		word[15'd6329] <= 32'd5405;
		word[15'd6330] <= 32'd5406;
		word[15'd6331] <= 32'd5407;
		word[15'd6332] <= 32'd5408;
		word[15'd6333] <= 32'd5409;
		word[15'd6334] <= 32'd5410;
		word[15'd6335] <= 32'd5411;
		word[15'd6336] <= 32'd5412;
		word[15'd6337] <= 32'd5413;
		word[15'd6338] <= 32'd5414;
		word[15'd6339] <= 32'd5415;
		word[15'd6340] <= 32'd5416;
		word[15'd6341] <= 32'd5417;
		word[15'd6342] <= 32'd5418;
		word[15'd6343] <= 32'd5419;
		word[15'd6344] <= 32'd5420;
		word[15'd6345] <= 32'd5421;
		word[15'd6346] <= 32'd5422;
		word[15'd6347] <= 32'd5423;
		word[15'd6348] <= 32'd5424;
		word[15'd6349] <= 32'd5425;
		word[15'd6350] <= 32'd5426;
		word[15'd6351] <= 32'd5427;
		word[15'd6352] <= 32'd5428;
		word[15'd6353] <= 32'd5429;
		word[15'd6354] <= 32'd5430;
		word[15'd6355] <= 32'd5431;
		word[15'd6356] <= 32'd5432;
		word[15'd6357] <= 32'd5433;
		word[15'd6358] <= 32'd5434;
		word[15'd6359] <= 32'd5435;
		word[15'd6360] <= 32'd5436;
		word[15'd6361] <= 32'd5437;
		word[15'd6362] <= 32'd5438;
		word[15'd6363] <= 32'd5439;
		word[15'd6364] <= 32'd5440;
		word[15'd6365] <= 32'd5441;
		word[15'd6366] <= 32'd5442;
		word[15'd6367] <= 32'd5443;
		word[15'd6368] <= 32'd5444;
		word[15'd6369] <= 32'd5445;
		word[15'd6370] <= 32'd5446;
		word[15'd6371] <= 32'd5447;
		word[15'd6372] <= 32'd5448;
		word[15'd6373] <= 32'd5449;
		word[15'd6374] <= 32'd5450;
		word[15'd6375] <= 32'd5451;
		word[15'd6376] <= 32'd5452;
		word[15'd6377] <= 32'd5453;
		word[15'd6378] <= 32'd5454;
		word[15'd6379] <= 32'd5455;
		word[15'd6380] <= 32'd5456;
		word[15'd6381] <= 32'd5457;
		word[15'd6382] <= 32'd5458;
		word[15'd6383] <= 32'd5459;
		word[15'd6384] <= 32'd5460;
		word[15'd6385] <= 32'd5461;
		word[15'd6386] <= 32'd5462;
		word[15'd6387] <= 32'd5463;
		word[15'd6388] <= 32'd5464;
		word[15'd6389] <= 32'd5465;
		word[15'd6390] <= 32'd5466;
		word[15'd6391] <= 32'd5467;
		word[15'd6392] <= 32'd5468;
		word[15'd6393] <= 32'd5469;
		word[15'd6394] <= 32'd5470;
		word[15'd6395] <= 32'd5471;
		word[15'd6396] <= 32'd5472;
		word[15'd6397] <= 32'd5473;
		word[15'd6398] <= 32'd5474;
		word[15'd6399] <= 32'd5475;
		word[15'd6400] <= 32'd5476;
		word[15'd6401] <= 32'd5477;
		word[15'd6402] <= 32'd5478;
		word[15'd6403] <= 32'd5479;
		word[15'd6404] <= 32'd5480;
		word[15'd6405] <= 32'd5481;
		word[15'd6406] <= 32'd5482;
		word[15'd6407] <= 32'd5483;
		word[15'd6408] <= 32'd5484;
		word[15'd6409] <= 32'd5485;
		word[15'd6410] <= 32'd5486;
		word[15'd6411] <= 32'd5487;
		word[15'd6412] <= 32'd5488;
		word[15'd6413] <= 32'd5489;
		word[15'd6414] <= 32'd5490;
		word[15'd6415] <= 32'd5491;
		word[15'd6416] <= 32'd5492;
		word[15'd6417] <= 32'd5493;
		word[15'd6418] <= 32'd5494;
		word[15'd6419] <= 32'd5495;
		word[15'd6420] <= 32'd5496;
		word[15'd6421] <= 32'd5497;
		word[15'd6422] <= 32'd5498;
		word[15'd6423] <= 32'd5499;
		word[15'd6424] <= 32'd5500;
		word[15'd6425] <= 32'd5501;
		word[15'd6426] <= 32'd5502;
		word[15'd6427] <= 32'd5503;
		word[15'd6428] <= 32'd5504;
		word[15'd6429] <= 32'd5505;
		word[15'd6430] <= 32'd5506;
		word[15'd6431] <= 32'd5507;
		word[15'd6432] <= 32'd5508;
		word[15'd6433] <= 32'd5509;
		word[15'd6434] <= 32'd5510;
		word[15'd6435] <= 32'd5511;
		word[15'd6436] <= 32'd5512;
		word[15'd6437] <= 32'd5513;
		word[15'd6438] <= 32'd5514;
		word[15'd6439] <= 32'd5515;
		word[15'd6440] <= 32'd5516;
		word[15'd6441] <= 32'd5517;
		word[15'd6442] <= 32'd5518;
		word[15'd6443] <= 32'd5519;
		word[15'd6444] <= 32'd5520;
		word[15'd6445] <= 32'd5521;
		word[15'd6446] <= 32'd5522;
		word[15'd6447] <= 32'd5523;
		word[15'd6448] <= 32'd5524;
		word[15'd6449] <= 32'd5525;
		word[15'd6450] <= 32'd5526;
		word[15'd6451] <= 32'd5527;
		word[15'd6452] <= 32'd5528;
		word[15'd6453] <= 32'd5529;
		word[15'd6454] <= 32'd5530;
		word[15'd6455] <= 32'd5531;
		word[15'd6456] <= 32'd5532;
		word[15'd6457] <= 32'd5533;
		word[15'd6458] <= 32'd5534;
		word[15'd6459] <= 32'd5535;
		word[15'd6460] <= 32'd5536;
		word[15'd6461] <= 32'd5537;
		word[15'd6462] <= 32'd5538;
		word[15'd6463] <= 32'd5539;
		word[15'd6464] <= 32'd5540;
		word[15'd6465] <= 32'd5541;
		word[15'd6466] <= 32'd5542;
		word[15'd6467] <= 32'd5543;
		word[15'd6468] <= 32'd5544;
		word[15'd6469] <= 32'd5545;
		word[15'd6470] <= 32'd5546;
		word[15'd6471] <= 32'd5547;
		word[15'd6472] <= 32'd5548;
		word[15'd6473] <= 32'd5549;
		word[15'd6474] <= 32'd5550;
		word[15'd6475] <= 32'd5551;
		word[15'd6476] <= 32'd5552;
		word[15'd6477] <= 32'd5553;
		word[15'd6478] <= 32'd5554;
		word[15'd6479] <= 32'd5555;
		word[15'd6480] <= 32'd5556;
		word[15'd6481] <= 32'd5557;
		word[15'd6482] <= 32'd5558;
		word[15'd6483] <= 32'd5559;
		word[15'd6484] <= 32'd5560;
		word[15'd6485] <= 32'd5561;
		word[15'd6486] <= 32'd5562;
		word[15'd6487] <= 32'd5563;
		word[15'd6488] <= 32'd5564;
		word[15'd6489] <= 32'd5565;
		word[15'd6490] <= 32'd5566;
		word[15'd6491] <= 32'd5567;
		word[15'd6492] <= 32'd5568;
		word[15'd6493] <= 32'd5569;
		word[15'd6494] <= 32'd5570;
		word[15'd6495] <= 32'd5571;
		word[15'd6496] <= 32'd5572;
		word[15'd6497] <= 32'd5573;
		word[15'd6498] <= 32'd5574;
		word[15'd6499] <= 32'd5575;
		word[15'd6500] <= 32'd5576;
		word[15'd6501] <= 32'd5577;
		word[15'd6502] <= 32'd5578;
		word[15'd6503] <= 32'd5579;
		word[15'd6504] <= 32'd5580;
		word[15'd6505] <= 32'd5581;
		word[15'd6506] <= 32'd5582;
		word[15'd6507] <= 32'd5583;
		word[15'd6508] <= 32'd5584;
		word[15'd6509] <= 32'd5585;
		word[15'd6510] <= 32'd5586;
		word[15'd6511] <= 32'd5587;
		word[15'd6512] <= 32'd5588;
		word[15'd6513] <= 32'd5589;
		word[15'd6514] <= 32'd5590;
		word[15'd6515] <= 32'd5591;
		word[15'd6516] <= 32'd5592;
		word[15'd6517] <= 32'd5593;
		word[15'd6518] <= 32'd5594;
		word[15'd6519] <= 32'd5595;
		word[15'd6520] <= 32'd5596;
		word[15'd6521] <= 32'd5597;
		word[15'd6522] <= 32'd5598;
		word[15'd6523] <= 32'd5599;
		word[15'd6524] <= 32'd5600;
		word[15'd6525] <= 32'd5601;
		word[15'd6526] <= 32'd5602;
		word[15'd6527] <= 32'd5603;
		word[15'd6528] <= 32'd5604;
		word[15'd6529] <= 32'd5605;
		word[15'd6530] <= 32'd5606;
		word[15'd6531] <= 32'd5607;
		word[15'd6532] <= 32'd5608;
		word[15'd6533] <= 32'd5609;
		word[15'd6534] <= 32'd5610;
		word[15'd6535] <= 32'd5611;
		word[15'd6536] <= 32'd5612;
		word[15'd6537] <= 32'd5613;
		word[15'd6538] <= 32'd5614;
		word[15'd6539] <= 32'd5615;
		word[15'd6540] <= 32'd5616;
		word[15'd6541] <= 32'd5617;
		word[15'd6542] <= 32'd5618;
		word[15'd6543] <= 32'd5619;
		word[15'd6544] <= 32'd5620;
		word[15'd6545] <= 32'd5621;
		word[15'd6546] <= 32'd5622;
		word[15'd6547] <= 32'd5623;
		word[15'd6548] <= 32'd5624;
		word[15'd6549] <= 32'd5625;
		word[15'd6550] <= 32'd5626;
		word[15'd6551] <= 32'd5627;
		word[15'd6552] <= 32'd5628;
		word[15'd6553] <= 32'd5629;
		word[15'd6554] <= 32'd5630;
		word[15'd6555] <= 32'd5631;
		word[15'd6556] <= 32'd5632;
		word[15'd6557] <= 32'd5633;
		word[15'd6558] <= 32'd5634;
		word[15'd6559] <= 32'd5635;
		word[15'd6560] <= 32'd5636;
		word[15'd6561] <= 32'd5637;
		word[15'd6562] <= 32'd5638;
		word[15'd6563] <= 32'd5639;
		word[15'd6564] <= 32'd5640;
		word[15'd6565] <= 32'd5641;
		word[15'd6566] <= 32'd5642;
		word[15'd6567] <= 32'd5643;
		word[15'd6568] <= 32'd5644;
		word[15'd6569] <= 32'd5645;
		word[15'd6570] <= 32'd5646;
		word[15'd6571] <= 32'd5647;
		word[15'd6572] <= 32'd5648;
		word[15'd6573] <= 32'd5649;
		word[15'd6574] <= 32'd5650;
		word[15'd6575] <= 32'd5651;
		word[15'd6576] <= 32'd5652;
		word[15'd6577] <= 32'd5653;
		word[15'd6578] <= 32'd5654;
		word[15'd6579] <= 32'd5655;
		word[15'd6580] <= 32'd5656;
		word[15'd6581] <= 32'd5657;
		word[15'd6582] <= 32'd5658;
		word[15'd6583] <= 32'd5659;
		word[15'd6584] <= 32'd5660;
		word[15'd6585] <= 32'd5661;
		word[15'd6586] <= 32'd5662;
		word[15'd6587] <= 32'd5663;
		word[15'd6588] <= 32'd5664;
		word[15'd6589] <= 32'd5665;
		word[15'd6590] <= 32'd5666;
		word[15'd6591] <= 32'd5667;
		word[15'd6592] <= 32'd5668;
		word[15'd6593] <= 32'd5669;
		word[15'd6594] <= 32'd5670;
		word[15'd6595] <= 32'd5671;
		word[15'd6596] <= 32'd5672;
		word[15'd6597] <= 32'd5673;
		word[15'd6598] <= 32'd5674;
		word[15'd6599] <= 32'd5675;
		word[15'd6600] <= 32'd5676;
		word[15'd6601] <= 32'd5677;
		word[15'd6602] <= 32'd5678;
		word[15'd6603] <= 32'd5679;
		word[15'd6604] <= 32'd5680;
		word[15'd6605] <= 32'd5681;
		word[15'd6606] <= 32'd5682;
		word[15'd6607] <= 32'd5683;
		word[15'd6608] <= 32'd5684;
		word[15'd6609] <= 32'd5685;
		word[15'd6610] <= 32'd5686;
		word[15'd6611] <= 32'd5687;
		word[15'd6612] <= 32'd5688;
		word[15'd6613] <= 32'd5689;
		word[15'd6614] <= 32'd5690;
		word[15'd6615] <= 32'd5691;
		word[15'd6616] <= 32'd5692;
		word[15'd6617] <= 32'd5693;
		word[15'd6618] <= 32'd5694;
		word[15'd6619] <= 32'd5695;
		word[15'd6620] <= 32'd5696;
		word[15'd6621] <= 32'd5697;
		word[15'd6622] <= 32'd5698;
		word[15'd6623] <= 32'd5699;
		word[15'd6624] <= 32'd5700;
		word[15'd6625] <= 32'd5701;
		word[15'd6626] <= 32'd5702;
		word[15'd6627] <= 32'd5703;
		word[15'd6628] <= 32'd5704;
		word[15'd6629] <= 32'd5705;
		word[15'd6630] <= 32'd5706;
		word[15'd6631] <= 32'd5707;
		word[15'd6632] <= 32'd5708;
		word[15'd6633] <= 32'd5709;
		word[15'd6634] <= 32'd5710;
		word[15'd6635] <= 32'd5711;
		word[15'd6636] <= 32'd5712;
		word[15'd6637] <= 32'd5713;
		word[15'd6638] <= 32'd5714;
		word[15'd6639] <= 32'd5715;
		word[15'd6640] <= 32'd5716;
		word[15'd6641] <= 32'd5717;
		word[15'd6642] <= 32'd5718;
		word[15'd6643] <= 32'd5719;
		word[15'd6644] <= 32'd5720;
		word[15'd6645] <= 32'd5721;
		word[15'd6646] <= 32'd5722;
		word[15'd6647] <= 32'd5723;
		word[15'd6648] <= 32'd5724;
		word[15'd6649] <= 32'd5725;
		word[15'd6650] <= 32'd5726;
		word[15'd6651] <= 32'd5727;
		word[15'd6652] <= 32'd5728;
		word[15'd6653] <= 32'd5729;
		word[15'd6654] <= 32'd5730;
		word[15'd6655] <= 32'd5731;
		word[15'd6656] <= 32'd5732;
		word[15'd6657] <= 32'd5733;
		word[15'd6658] <= 32'd5734;
		word[15'd6659] <= 32'd5735;
		word[15'd6660] <= 32'd5736;
		word[15'd6661] <= 32'd5737;
		word[15'd6662] <= 32'd5738;
		word[15'd6663] <= 32'd5739;
		word[15'd6664] <= 32'd5740;
		word[15'd6665] <= 32'd5741;
		word[15'd6666] <= 32'd5742;
		word[15'd6667] <= 32'd5743;
		word[15'd6668] <= 32'd5744;
		word[15'd6669] <= 32'd5745;
		word[15'd6670] <= 32'd5746;
		word[15'd6671] <= 32'd5747;
		word[15'd6672] <= 32'd5748;
		word[15'd6673] <= 32'd5749;
		word[15'd6674] <= 32'd5750;
		word[15'd6675] <= 32'd5751;
		word[15'd6676] <= 32'd5752;
		word[15'd6677] <= 32'd5753;
		word[15'd6678] <= 32'd5754;
		word[15'd6679] <= 32'd5755;
		word[15'd6680] <= 32'd5756;
		word[15'd6681] <= 32'd5757;
		word[15'd6682] <= 32'd5758;
		word[15'd6683] <= 32'd5759;
		word[15'd6684] <= 32'd5760;
		word[15'd6685] <= 32'd5761;
		word[15'd6686] <= 32'd5762;
		word[15'd6687] <= 32'd5763;
		word[15'd6688] <= 32'd5764;
		word[15'd6689] <= 32'd5765;
		word[15'd6690] <= 32'd5766;
		word[15'd6691] <= 32'd5767;
		word[15'd6692] <= 32'd5768;
		word[15'd6693] <= 32'd5769;
		word[15'd6694] <= 32'd5770;
		word[15'd6695] <= 32'd5771;
		word[15'd6696] <= 32'd5772;
		word[15'd6697] <= 32'd5773;
		word[15'd6698] <= 32'd5774;
		word[15'd6699] <= 32'd5775;
		word[15'd6700] <= 32'd5776;
		word[15'd6701] <= 32'd5777;
		word[15'd6702] <= 32'd5778;
		word[15'd6703] <= 32'd5779;
		word[15'd6704] <= 32'd5780;
		word[15'd6705] <= 32'd5781;
		word[15'd6706] <= 32'd5782;
		word[15'd6707] <= 32'd5783;
		word[15'd6708] <= 32'd5784;
		word[15'd6709] <= 32'd5785;
		word[15'd6710] <= 32'd5786;
		word[15'd6711] <= 32'd5787;
		word[15'd6712] <= 32'd5788;
		word[15'd6713] <= 32'd5789;
		word[15'd6714] <= 32'd5790;
		word[15'd6715] <= 32'd5791;
		word[15'd6716] <= 32'd5792;
		word[15'd6717] <= 32'd5793;
		word[15'd6718] <= 32'd5794;
		word[15'd6719] <= 32'd5795;
		word[15'd6720] <= 32'd5796;
		word[15'd6721] <= 32'd5797;
		word[15'd6722] <= 32'd5798;
		word[15'd6723] <= 32'd5799;
		word[15'd6724] <= 32'd5800;
		word[15'd6725] <= 32'd5801;
		word[15'd6726] <= 32'd5802;
		word[15'd6727] <= 32'd5803;
		word[15'd6728] <= 32'd5804;
		word[15'd6729] <= 32'd5805;
		word[15'd6730] <= 32'd5806;
		word[15'd6731] <= 32'd5807;
		word[15'd6732] <= 32'd5808;
		word[15'd6733] <= 32'd5809;
		word[15'd6734] <= 32'd5810;
		word[15'd6735] <= 32'd5811;
		word[15'd6736] <= 32'd5812;
		word[15'd6737] <= 32'd5813;
		word[15'd6738] <= 32'd5814;
		word[15'd6739] <= 32'd5815;
		word[15'd6740] <= 32'd5816;
		word[15'd6741] <= 32'd5817;
		word[15'd6742] <= 32'd5818;
		word[15'd6743] <= 32'd5819;
		word[15'd6744] <= 32'd5820;
		word[15'd6745] <= 32'd5821;
		word[15'd6746] <= 32'd5822;
		word[15'd6747] <= 32'd5823;
		word[15'd6748] <= 32'd5824;
		word[15'd6749] <= 32'd5825;
		word[15'd6750] <= 32'd5826;
		word[15'd6751] <= 32'd5827;
		word[15'd6752] <= 32'd5828;
		word[15'd6753] <= 32'd5829;
		word[15'd6754] <= 32'd5830;
		word[15'd6755] <= 32'd5831;
		word[15'd6756] <= 32'd5832;
		word[15'd6757] <= 32'd5833;
		word[15'd6758] <= 32'd5834;
		word[15'd6759] <= 32'd5835;
		word[15'd6760] <= 32'd5836;
		word[15'd6761] <= 32'd5837;
		word[15'd6762] <= 32'd5838;
		word[15'd6763] <= 32'd5839;
		word[15'd6764] <= 32'd5840;
		word[15'd6765] <= 32'd5841;
		word[15'd6766] <= 32'd5842;
		word[15'd6767] <= 32'd5843;
		word[15'd6768] <= 32'd5844;
		word[15'd6769] <= 32'd5845;
		word[15'd6770] <= 32'd5846;
		word[15'd6771] <= 32'd5847;
		word[15'd6772] <= 32'd5848;
		word[15'd6773] <= 32'd5849;
		word[15'd6774] <= 32'd5850;
		word[15'd6775] <= 32'd5851;
		word[15'd6776] <= 32'd5852;
		word[15'd6777] <= 32'd5853;
		word[15'd6778] <= 32'd5854;
		word[15'd6779] <= 32'd5855;
		word[15'd6780] <= 32'd5856;
		word[15'd6781] <= 32'd5857;
		word[15'd6782] <= 32'd5858;
		word[15'd6783] <= 32'd5859;
		word[15'd6784] <= 32'd5860;
		word[15'd6785] <= 32'd5861;
		word[15'd6786] <= 32'd5862;
		word[15'd6787] <= 32'd5863;
		word[15'd6788] <= 32'd5864;
		word[15'd6789] <= 32'd5865;
		word[15'd6790] <= 32'd5866;
		word[15'd6791] <= 32'd5867;
		word[15'd6792] <= 32'd5868;
		word[15'd6793] <= 32'd5869;
		word[15'd6794] <= 32'd5870;
		word[15'd6795] <= 32'd5871;
		word[15'd6796] <= 32'd5872;
		word[15'd6797] <= 32'd5873;
		word[15'd6798] <= 32'd5874;
		word[15'd6799] <= 32'd5875;
		word[15'd6800] <= 32'd5876;
		word[15'd6801] <= 32'd5877;
		word[15'd6802] <= 32'd5878;
		word[15'd6803] <= 32'd5879;
		word[15'd6804] <= 32'd5880;
		word[15'd6805] <= 32'd5881;
		word[15'd6806] <= 32'd5882;
		word[15'd6807] <= 32'd5883;
		word[15'd6808] <= 32'd5884;
		word[15'd6809] <= 32'd5885;
		word[15'd6810] <= 32'd5886;
		word[15'd6811] <= 32'd5887;
		word[15'd6812] <= 32'd5888;
		word[15'd6813] <= 32'd5889;
		word[15'd6814] <= 32'd5890;
		word[15'd6815] <= 32'd5891;
		word[15'd6816] <= 32'd5892;
		word[15'd6817] <= 32'd5893;
		word[15'd6818] <= 32'd5894;
		word[15'd6819] <= 32'd5895;
		word[15'd6820] <= 32'd5896;
		word[15'd6821] <= 32'd5897;
		word[15'd6822] <= 32'd5898;
		word[15'd6823] <= 32'd5899;
		word[15'd6824] <= 32'd5900;
		word[15'd6825] <= 32'd5901;
		word[15'd6826] <= 32'd5902;
		word[15'd6827] <= 32'd5903;
		word[15'd6828] <= 32'd5904;
		word[15'd6829] <= 32'd5905;
		word[15'd6830] <= 32'd5906;
		word[15'd6831] <= 32'd5907;
		word[15'd6832] <= 32'd5908;
		word[15'd6833] <= 32'd5909;
		word[15'd6834] <= 32'd5910;
		word[15'd6835] <= 32'd5911;
		word[15'd6836] <= 32'd5912;
		word[15'd6837] <= 32'd5913;
		word[15'd6838] <= 32'd5914;
		word[15'd6839] <= 32'd5915;
		word[15'd6840] <= 32'd5916;
		word[15'd6841] <= 32'd5917;
		word[15'd6842] <= 32'd5918;
		word[15'd6843] <= 32'd5919;
		word[15'd6844] <= 32'd5920;
		word[15'd6845] <= 32'd5921;
		word[15'd6846] <= 32'd5922;
		word[15'd6847] <= 32'd5923;
		word[15'd6848] <= 32'd5924;
		word[15'd6849] <= 32'd5925;
		word[15'd6850] <= 32'd5926;
		word[15'd6851] <= 32'd5927;
		word[15'd6852] <= 32'd5928;
		word[15'd6853] <= 32'd5929;
		word[15'd6854] <= 32'd5930;
		word[15'd6855] <= 32'd5931;
		word[15'd6856] <= 32'd5932;
		word[15'd6857] <= 32'd5933;
		word[15'd6858] <= 32'd5934;
		word[15'd6859] <= 32'd5935;
		word[15'd6860] <= 32'd5936;
		word[15'd6861] <= 32'd5937;
		word[15'd6862] <= 32'd5938;
		word[15'd6863] <= 32'd5939;
		word[15'd6864] <= 32'd5940;
		word[15'd6865] <= 32'd5941;
		word[15'd6866] <= 32'd5942;
		word[15'd6867] <= 32'd5943;
		word[15'd6868] <= 32'd5944;
		word[15'd6869] <= 32'd5945;
		word[15'd6870] <= 32'd5946;
		word[15'd6871] <= 32'd5947;
		word[15'd6872] <= 32'd5948;
		word[15'd6873] <= 32'd5949;
		word[15'd6874] <= 32'd5950;
		word[15'd6875] <= 32'd5951;
		word[15'd6876] <= 32'd5952;
		word[15'd6877] <= 32'd5953;
		word[15'd6878] <= 32'd5954;
		word[15'd6879] <= 32'd5955;
		word[15'd6880] <= 32'd5956;
		word[15'd6881] <= 32'd5957;
		word[15'd6882] <= 32'd5958;
		word[15'd6883] <= 32'd5959;
		word[15'd6884] <= 32'd5960;
		word[15'd6885] <= 32'd5961;
		word[15'd6886] <= 32'd5962;
		word[15'd6887] <= 32'd5963;
		word[15'd6888] <= 32'd5964;
		word[15'd6889] <= 32'd5965;
		word[15'd6890] <= 32'd5966;
		word[15'd6891] <= 32'd5967;
		word[15'd6892] <= 32'd5968;
		word[15'd6893] <= 32'd5969;
		word[15'd6894] <= 32'd5970;
		word[15'd6895] <= 32'd5971;
		word[15'd6896] <= 32'd5972;
		word[15'd6897] <= 32'd5973;
		word[15'd6898] <= 32'd5974;
		word[15'd6899] <= 32'd5975;
		word[15'd6900] <= 32'd5976;
		word[15'd6901] <= 32'd5977;
		word[15'd6902] <= 32'd5978;
		word[15'd6903] <= 32'd5979;
		word[15'd6904] <= 32'd5980;
		word[15'd6905] <= 32'd5981;
		word[15'd6906] <= 32'd5982;
		word[15'd6907] <= 32'd5983;
		word[15'd6908] <= 32'd5984;
		word[15'd6909] <= 32'd5985;
		word[15'd6910] <= 32'd5986;
		word[15'd6911] <= 32'd5987;
		word[15'd6912] <= 32'd5988;
		word[15'd6913] <= 32'd5989;
		word[15'd6914] <= 32'd5990;
		word[15'd6915] <= 32'd5991;
		word[15'd6916] <= 32'd5992;
		word[15'd6917] <= 32'd5993;
		word[15'd6918] <= 32'd5994;
		word[15'd6919] <= 32'd5995;
		word[15'd6920] <= 32'd5996;
		word[15'd6921] <= 32'd5997;
		word[15'd6922] <= 32'd5998;
		word[15'd6923] <= 32'd5999;
		word[15'd6924] <= 32'd6000;
		word[15'd6925] <= 32'd6001;
		word[15'd6926] <= 32'd6002;
		word[15'd6927] <= 32'd6003;
		word[15'd6928] <= 32'd6004;
		word[15'd6929] <= 32'd6005;
		word[15'd6930] <= 32'd6006;
		word[15'd6931] <= 32'd6007;
		word[15'd6932] <= 32'd6008;
		word[15'd6933] <= 32'd6009;
		word[15'd6934] <= 32'd6010;
		word[15'd6935] <= 32'd6011;
		word[15'd6936] <= 32'd6012;
		word[15'd6937] <= 32'd6013;
		word[15'd6938] <= 32'd6014;
		word[15'd6939] <= 32'd6015;
		word[15'd6940] <= 32'd6016;
		word[15'd6941] <= 32'd6017;
		word[15'd6942] <= 32'd6018;
		word[15'd6943] <= 32'd6019;
		word[15'd6944] <= 32'd6020;
		word[15'd6945] <= 32'd6021;
		word[15'd6946] <= 32'd6022;
		word[15'd6947] <= 32'd6023;
		word[15'd6948] <= 32'd6024;
		word[15'd6949] <= 32'd6025;
		word[15'd6950] <= 32'd6026;
		word[15'd6951] <= 32'd6027;
		word[15'd6952] <= 32'd6028;
		word[15'd6953] <= 32'd6029;
		word[15'd6954] <= 32'd6030;
		word[15'd6955] <= 32'd6031;
		word[15'd6956] <= 32'd6032;
		word[15'd6957] <= 32'd6033;
		word[15'd6958] <= 32'd6034;
		word[15'd6959] <= 32'd6035;
		word[15'd6960] <= 32'd6036;
		word[15'd6961] <= 32'd6037;
		word[15'd6962] <= 32'd6038;
		word[15'd6963] <= 32'd6039;
		word[15'd6964] <= 32'd6040;
		word[15'd6965] <= 32'd6041;
		word[15'd6966] <= 32'd6042;
		word[15'd6967] <= 32'd6043;
		word[15'd6968] <= 32'd6044;
		word[15'd6969] <= 32'd6045;
		word[15'd6970] <= 32'd6046;
		word[15'd6971] <= 32'd6047;
		word[15'd6972] <= 32'd6048;
		word[15'd6973] <= 32'd6049;
		word[15'd6974] <= 32'd6050;
		word[15'd6975] <= 32'd6051;
		word[15'd6976] <= 32'd6052;
		word[15'd6977] <= 32'd6053;
		word[15'd6978] <= 32'd6054;
		word[15'd6979] <= 32'd6055;
		word[15'd6980] <= 32'd6056;
		word[15'd6981] <= 32'd6057;
		word[15'd6982] <= 32'd6058;
		word[15'd6983] <= 32'd6059;
		word[15'd6984] <= 32'd6060;
		word[15'd6985] <= 32'd6061;
		word[15'd6986] <= 32'd6062;
		word[15'd6987] <= 32'd6063;
		word[15'd6988] <= 32'd6064;
		word[15'd6989] <= 32'd6065;
		word[15'd6990] <= 32'd6066;
		word[15'd6991] <= 32'd6067;
		word[15'd6992] <= 32'd6068;
		word[15'd6993] <= 32'd6069;
		word[15'd6994] <= 32'd6070;
		word[15'd6995] <= 32'd6071;
		word[15'd6996] <= 32'd6072;
		word[15'd6997] <= 32'd6073;
		word[15'd6998] <= 32'd6074;
		word[15'd6999] <= 32'd6075;
		word[15'd7000] <= 32'd6076;
		word[15'd7001] <= 32'd6077;
		word[15'd7002] <= 32'd6078;
		word[15'd7003] <= 32'd6079;
		word[15'd7004] <= 32'd6080;
		word[15'd7005] <= 32'd6081;
		word[15'd7006] <= 32'd6082;
		word[15'd7007] <= 32'd6083;
		word[15'd7008] <= 32'd6084;
		word[15'd7009] <= 32'd6085;
		word[15'd7010] <= 32'd6086;
		word[15'd7011] <= 32'd6087;
		word[15'd7012] <= 32'd6088;
		word[15'd7013] <= 32'd6089;
		word[15'd7014] <= 32'd6090;
		word[15'd7015] <= 32'd6091;
		word[15'd7016] <= 32'd6092;
		word[15'd7017] <= 32'd6093;
		word[15'd7018] <= 32'd6094;
		word[15'd7019] <= 32'd6095;
		word[15'd7020] <= 32'd6096;
		word[15'd7021] <= 32'd6097;
		word[15'd7022] <= 32'd6098;
		word[15'd7023] <= 32'd6099;
		word[15'd7024] <= 32'd6100;
		word[15'd7025] <= 32'd6101;
		word[15'd7026] <= 32'd6102;
		word[15'd7027] <= 32'd6103;
		word[15'd7028] <= 32'd6104;
		word[15'd7029] <= 32'd6105;
		word[15'd7030] <= 32'd6106;
		word[15'd7031] <= 32'd6107;
		word[15'd7032] <= 32'd6108;
		word[15'd7033] <= 32'd6109;
		word[15'd7034] <= 32'd6110;
		word[15'd7035] <= 32'd6111;
		word[15'd7036] <= 32'd6112;
		word[15'd7037] <= 32'd6113;
		word[15'd7038] <= 32'd6114;
		word[15'd7039] <= 32'd6115;
		word[15'd7040] <= 32'd6116;
		word[15'd7041] <= 32'd6117;
		word[15'd7042] <= 32'd6118;
		word[15'd7043] <= 32'd6119;
		word[15'd7044] <= 32'd6120;
		word[15'd7045] <= 32'd6121;
		word[15'd7046] <= 32'd6122;
		word[15'd7047] <= 32'd6123;
		word[15'd7048] <= 32'd6124;
		word[15'd7049] <= 32'd6125;
		word[15'd7050] <= 32'd6126;
		word[15'd7051] <= 32'd6127;
		word[15'd7052] <= 32'd6128;
		word[15'd7053] <= 32'd6129;
		word[15'd7054] <= 32'd6130;
		word[15'd7055] <= 32'd6131;
		word[15'd7056] <= 32'd6132;
		word[15'd7057] <= 32'd6133;
		word[15'd7058] <= 32'd6134;
		word[15'd7059] <= 32'd6135;
		word[15'd7060] <= 32'd6136;
		word[15'd7061] <= 32'd6137;
		word[15'd7062] <= 32'd6138;
		word[15'd7063] <= 32'd6139;
		word[15'd7064] <= 32'd6140;
		word[15'd7065] <= 32'd6141;
		word[15'd7066] <= 32'd6142;
		word[15'd7067] <= 32'd6143;
		word[15'd7068] <= 32'd6144;
		word[15'd7069] <= 32'd6145;
		word[15'd7070] <= 32'd6146;
		word[15'd7071] <= 32'd6147;
		word[15'd7072] <= 32'd6148;
		word[15'd7073] <= 32'd6149;
		word[15'd7074] <= 32'd6150;
		word[15'd7075] <= 32'd6151;
		word[15'd7076] <= 32'd6152;
		word[15'd7077] <= 32'd6153;
		word[15'd7078] <= 32'd6154;
		word[15'd7079] <= 32'd6155;
		word[15'd7080] <= 32'd6156;
		word[15'd7081] <= 32'd6157;
		word[15'd7082] <= 32'd6158;
		word[15'd7083] <= 32'd6159;
		word[15'd7084] <= 32'd6160;
		word[15'd7085] <= 32'd6161;
		word[15'd7086] <= 32'd6162;
		word[15'd7087] <= 32'd6163;
		word[15'd7088] <= 32'd6164;
		word[15'd7089] <= 32'd6165;
		word[15'd7090] <= 32'd6166;
		word[15'd7091] <= 32'd6167;
		word[15'd7092] <= 32'd6168;
		word[15'd7093] <= 32'd6169;
		word[15'd7094] <= 32'd6170;
		word[15'd7095] <= 32'd6171;
		word[15'd7096] <= 32'd6172;
		word[15'd7097] <= 32'd6173;
		word[15'd7098] <= 32'd6174;
		word[15'd7099] <= 32'd6175;
		word[15'd7100] <= 32'd6176;
		word[15'd7101] <= 32'd6177;
		word[15'd7102] <= 32'd6178;
		word[15'd7103] <= 32'd6179;
		word[15'd7104] <= 32'd6180;
		word[15'd7105] <= 32'd6181;
		word[15'd7106] <= 32'd6182;
		word[15'd7107] <= 32'd6183;
		word[15'd7108] <= 32'd6184;
		word[15'd7109] <= 32'd6185;
		word[15'd7110] <= 32'd6186;
		word[15'd7111] <= 32'd6187;
		word[15'd7112] <= 32'd6188;
		word[15'd7113] <= 32'd6189;
		word[15'd7114] <= 32'd6190;
		word[15'd7115] <= 32'd6191;
		word[15'd7116] <= 32'd6192;
		word[15'd7117] <= 32'd6193;
		word[15'd7118] <= 32'd6194;
		word[15'd7119] <= 32'd6195;
		word[15'd7120] <= 32'd6196;
		word[15'd7121] <= 32'd6197;
		word[15'd7122] <= 32'd6198;
		word[15'd7123] <= 32'd6199;
		word[15'd7124] <= 32'd6200;
		word[15'd7125] <= 32'd6201;
		word[15'd7126] <= 32'd6202;
		word[15'd7127] <= 32'd6203;
		word[15'd7128] <= 32'd6204;
		word[15'd7129] <= 32'd6205;
		word[15'd7130] <= 32'd6206;
		word[15'd7131] <= 32'd6207;
		word[15'd7132] <= 32'd6208;
		word[15'd7133] <= 32'd6209;
		word[15'd7134] <= 32'd6210;
		word[15'd7135] <= 32'd6211;
		word[15'd7136] <= 32'd6212;
		word[15'd7137] <= 32'd6213;
		word[15'd7138] <= 32'd6214;
		word[15'd7139] <= 32'd6215;
		word[15'd7140] <= 32'd6216;
		word[15'd7141] <= 32'd6217;
		word[15'd7142] <= 32'd6218;
		word[15'd7143] <= 32'd6219;
		word[15'd7144] <= 32'd6220;
		word[15'd7145] <= 32'd6221;
		word[15'd7146] <= 32'd6222;
		word[15'd7147] <= 32'd6223;
		word[15'd7148] <= 32'd6224;
		word[15'd7149] <= 32'd6225;
		word[15'd7150] <= 32'd6226;
		word[15'd7151] <= 32'd6227;
		word[15'd7152] <= 32'd6228;
		word[15'd7153] <= 32'd6229;
		word[15'd7154] <= 32'd6230;
		word[15'd7155] <= 32'd6231;
		word[15'd7156] <= 32'd6232;
		word[15'd7157] <= 32'd6233;
		word[15'd7158] <= 32'd6234;
		word[15'd7159] <= 32'd6235;
		word[15'd7160] <= 32'd6236;
		word[15'd7161] <= 32'd6237;
		word[15'd7162] <= 32'd6238;
		word[15'd7163] <= 32'd6239;
		word[15'd7164] <= 32'd6240;
		word[15'd7165] <= 32'd6241;
		word[15'd7166] <= 32'd6242;
		word[15'd7167] <= 32'd6243;
		word[15'd7168] <= 32'd6244;
		word[15'd7169] <= 32'd6245;
		word[15'd7170] <= 32'd6246;
		word[15'd7171] <= 32'd6247;
		word[15'd7172] <= 32'd6248;
		word[15'd7173] <= 32'd6249;
		word[15'd7174] <= 32'd6250;
		word[15'd7175] <= 32'd6251;
		word[15'd7176] <= 32'd6252;
		word[15'd7177] <= 32'd6253;
		word[15'd7178] <= 32'd6254;
		word[15'd7179] <= 32'd6255;
		word[15'd7180] <= 32'd6256;
		word[15'd7181] <= 32'd6257;
		word[15'd7182] <= 32'd6258;
		word[15'd7183] <= 32'd6259;
		word[15'd7184] <= 32'd6260;
		word[15'd7185] <= 32'd6261;
		word[15'd7186] <= 32'd6262;
		word[15'd7187] <= 32'd6263;
		word[15'd7188] <= 32'd6264;
		word[15'd7189] <= 32'd6265;
		word[15'd7190] <= 32'd6266;
		word[15'd7191] <= 32'd6267;
		word[15'd7192] <= 32'd6268;
		word[15'd7193] <= 32'd6269;
		word[15'd7194] <= 32'd6270;
		word[15'd7195] <= 32'd6271;
		word[15'd7196] <= 32'd6272;
		word[15'd7197] <= 32'd6273;
		word[15'd7198] <= 32'd6274;
		word[15'd7199] <= 32'd6275;
		word[15'd7200] <= 32'd6276;
		word[15'd7201] <= 32'd6277;
		word[15'd7202] <= 32'd6278;
		word[15'd7203] <= 32'd6279;
		word[15'd7204] <= 32'd6280;
		word[15'd7205] <= 32'd6281;
		word[15'd7206] <= 32'd6282;
		word[15'd7207] <= 32'd6283;
		word[15'd7208] <= 32'd6284;
		word[15'd7209] <= 32'd6285;
		word[15'd7210] <= 32'd6286;
		word[15'd7211] <= 32'd6287;
		word[15'd7212] <= 32'd6288;
		word[15'd7213] <= 32'd6289;
		word[15'd7214] <= 32'd6290;
		word[15'd7215] <= 32'd6291;
		word[15'd7216] <= 32'd6292;
		word[15'd7217] <= 32'd6293;
		word[15'd7218] <= 32'd6294;
		word[15'd7219] <= 32'd6295;
		word[15'd7220] <= 32'd6296;
		word[15'd7221] <= 32'd6297;
		word[15'd7222] <= 32'd6298;
		word[15'd7223] <= 32'd6299;
		word[15'd7224] <= 32'd6300;
		word[15'd7225] <= 32'd6301;
		word[15'd7226] <= 32'd6302;
		word[15'd7227] <= 32'd6303;
		word[15'd7228] <= 32'd6304;
		word[15'd7229] <= 32'd6305;
		word[15'd7230] <= 32'd6306;
		word[15'd7231] <= 32'd6307;
		word[15'd7232] <= 32'd6308;
		word[15'd7233] <= 32'd6309;
		word[15'd7234] <= 32'd6310;
		word[15'd7235] <= 32'd6311;
		word[15'd7236] <= 32'd6312;
		word[15'd7237] <= 32'd6313;
		word[15'd7238] <= 32'd6314;
		word[15'd7239] <= 32'd6315;
		word[15'd7240] <= 32'd6316;
		word[15'd7241] <= 32'd6317;
		word[15'd7242] <= 32'd6318;
		word[15'd7243] <= 32'd6319;
		word[15'd7244] <= 32'd6320;
		word[15'd7245] <= 32'd6321;
		word[15'd7246] <= 32'd6322;
		word[15'd7247] <= 32'd6323;
		word[15'd7248] <= 32'd6324;
		word[15'd7249] <= 32'd6325;
		word[15'd7250] <= 32'd6326;
		word[15'd7251] <= 32'd6327;
		word[15'd7252] <= 32'd6328;
		word[15'd7253] <= 32'd6329;
		word[15'd7254] <= 32'd6330;
		word[15'd7255] <= 32'd6331;
		word[15'd7256] <= 32'd6332;
		word[15'd7257] <= 32'd6333;
		word[15'd7258] <= 32'd6334;
		word[15'd7259] <= 32'd6335;
		word[15'd7260] <= 32'd6336;
		word[15'd7261] <= 32'd6337;
		word[15'd7262] <= 32'd6338;
		word[15'd7263] <= 32'd6339;
		word[15'd7264] <= 32'd6340;
		word[15'd7265] <= 32'd6341;
		word[15'd7266] <= 32'd6342;
		word[15'd7267] <= 32'd6343;
		word[15'd7268] <= 32'd6344;
		word[15'd7269] <= 32'd6345;
		word[15'd7270] <= 32'd6346;
		word[15'd7271] <= 32'd6347;
		word[15'd7272] <= 32'd6348;
		word[15'd7273] <= 32'd6349;
		word[15'd7274] <= 32'd6350;
		word[15'd7275] <= 32'd6351;
		word[15'd7276] <= 32'd6352;
		word[15'd7277] <= 32'd6353;
		word[15'd7278] <= 32'd6354;
		word[15'd7279] <= 32'd6355;
		word[15'd7280] <= 32'd6356;
		word[15'd7281] <= 32'd6357;
		word[15'd7282] <= 32'd6358;
		word[15'd7283] <= 32'd6359;
		word[15'd7284] <= 32'd6360;
		word[15'd7285] <= 32'd6361;
		word[15'd7286] <= 32'd6362;
		word[15'd7287] <= 32'd6363;
		word[15'd7288] <= 32'd6364;
		word[15'd7289] <= 32'd6365;
		word[15'd7290] <= 32'd6366;
		word[15'd7291] <= 32'd6367;
		word[15'd7292] <= 32'd6368;
		word[15'd7293] <= 32'd6369;
		word[15'd7294] <= 32'd6370;
		word[15'd7295] <= 32'd6371;
		word[15'd7296] <= 32'd6372;
		word[15'd7297] <= 32'd6373;
		word[15'd7298] <= 32'd6374;
		word[15'd7299] <= 32'd6375;
		word[15'd7300] <= 32'd6376;
		word[15'd7301] <= 32'd6377;
		word[15'd7302] <= 32'd6378;
		word[15'd7303] <= 32'd6379;
		word[15'd7304] <= 32'd6380;
		word[15'd7305] <= 32'd6381;
		word[15'd7306] <= 32'd6382;
		word[15'd7307] <= 32'd6383;
		word[15'd7308] <= 32'd6384;
		word[15'd7309] <= 32'd6385;
		word[15'd7310] <= 32'd6386;
		word[15'd7311] <= 32'd6387;
		word[15'd7312] <= 32'd6388;
		word[15'd7313] <= 32'd6389;
		word[15'd7314] <= 32'd6390;
		word[15'd7315] <= 32'd6391;
		word[15'd7316] <= 32'd6392;
		word[15'd7317] <= 32'd6393;
		word[15'd7318] <= 32'd6394;
		word[15'd7319] <= 32'd6395;
		word[15'd7320] <= 32'd6396;
		word[15'd7321] <= 32'd6397;
		word[15'd7322] <= 32'd6398;
		word[15'd7323] <= 32'd6399;
		word[15'd7324] <= 32'd6400;
		word[15'd7325] <= 32'd6401;
		word[15'd7326] <= 32'd6402;
		word[15'd7327] <= 32'd6403;
		word[15'd7328] <= 32'd6404;
		word[15'd7329] <= 32'd6405;
		word[15'd7330] <= 32'd6406;
		word[15'd7331] <= 32'd6407;
		word[15'd7332] <= 32'd6408;
		word[15'd7333] <= 32'd6409;
		word[15'd7334] <= 32'd6410;
		word[15'd7335] <= 32'd6411;
		word[15'd7336] <= 32'd6412;
		word[15'd7337] <= 32'd6413;
		word[15'd7338] <= 32'd6414;
		word[15'd7339] <= 32'd6415;
		word[15'd7340] <= 32'd6416;
		word[15'd7341] <= 32'd6417;
		word[15'd7342] <= 32'd6418;
		word[15'd7343] <= 32'd6419;
		word[15'd7344] <= 32'd6420;
		word[15'd7345] <= 32'd6421;
		word[15'd7346] <= 32'd6422;
		word[15'd7347] <= 32'd6423;
		word[15'd7348] <= 32'd6424;
		word[15'd7349] <= 32'd6425;
		word[15'd7350] <= 32'd6426;
		word[15'd7351] <= 32'd6427;
		word[15'd7352] <= 32'd6428;
		word[15'd7353] <= 32'd6429;
		word[15'd7354] <= 32'd6430;
		word[15'd7355] <= 32'd6431;
		word[15'd7356] <= 32'd6432;
		word[15'd7357] <= 32'd6433;
		word[15'd7358] <= 32'd6434;
		word[15'd7359] <= 32'd6435;
		word[15'd7360] <= 32'd6436;
		word[15'd7361] <= 32'd6437;
		word[15'd7362] <= 32'd6438;
		word[15'd7363] <= 32'd6439;
		word[15'd7364] <= 32'd6440;
		word[15'd7365] <= 32'd6441;
		word[15'd7366] <= 32'd6442;
		word[15'd7367] <= 32'd6443;
		word[15'd7368] <= 32'd6444;
		word[15'd7369] <= 32'd6445;
		word[15'd7370] <= 32'd6446;
		word[15'd7371] <= 32'd6447;
		word[15'd7372] <= 32'd6448;
		word[15'd7373] <= 32'd6449;
		word[15'd7374] <= 32'd6450;
		word[15'd7375] <= 32'd6451;
		word[15'd7376] <= 32'd6452;
		word[15'd7377] <= 32'd6453;
		word[15'd7378] <= 32'd6454;
		word[15'd7379] <= 32'd6455;
		word[15'd7380] <= 32'd6456;
		word[15'd7381] <= 32'd6457;
		word[15'd7382] <= 32'd6458;
		word[15'd7383] <= 32'd6459;
		word[15'd7384] <= 32'd6460;
		word[15'd7385] <= 32'd6461;
		word[15'd7386] <= 32'd6462;
		word[15'd7387] <= 32'd6463;
		word[15'd7388] <= 32'd6464;
		word[15'd7389] <= 32'd6465;
		word[15'd7390] <= 32'd6466;
		word[15'd7391] <= 32'd6467;
		word[15'd7392] <= 32'd6468;
		word[15'd7393] <= 32'd6469;
		word[15'd7394] <= 32'd6470;
		word[15'd7395] <= 32'd6471;
		word[15'd7396] <= 32'd6472;
		word[15'd7397] <= 32'd6473;
		word[15'd7398] <= 32'd6474;
		word[15'd7399] <= 32'd6475;
		word[15'd7400] <= 32'd6476;
		word[15'd7401] <= 32'd6477;
		word[15'd7402] <= 32'd6478;
		word[15'd7403] <= 32'd6479;
		word[15'd7404] <= 32'd6480;
		word[15'd7405] <= 32'd6481;
		word[15'd7406] <= 32'd6482;
		word[15'd7407] <= 32'd6483;
		word[15'd7408] <= 32'd6484;
		word[15'd7409] <= 32'd6485;
		word[15'd7410] <= 32'd6486;
		word[15'd7411] <= 32'd6487;
		word[15'd7412] <= 32'd6488;
		word[15'd7413] <= 32'd6489;
		word[15'd7414] <= 32'd6490;
		word[15'd7415] <= 32'd6491;
		word[15'd7416] <= 32'd6492;
		word[15'd7417] <= 32'd6493;
		word[15'd7418] <= 32'd6494;
		word[15'd7419] <= 32'd6495;
		word[15'd7420] <= 32'd6496;
		word[15'd7421] <= 32'd6497;
		word[15'd7422] <= 32'd6498;
		word[15'd7423] <= 32'd6499;
		word[15'd7424] <= 32'd6500;
		word[15'd7425] <= 32'd6501;
		word[15'd7426] <= 32'd6502;
		word[15'd7427] <= 32'd6503;
		word[15'd7428] <= 32'd6504;
		word[15'd7429] <= 32'd6505;
		word[15'd7430] <= 32'd6506;
		word[15'd7431] <= 32'd6507;
		word[15'd7432] <= 32'd6508;
		word[15'd7433] <= 32'd6509;
		word[15'd7434] <= 32'd6510;
		word[15'd7435] <= 32'd6511;
		word[15'd7436] <= 32'd6512;
		word[15'd7437] <= 32'd6513;
		word[15'd7438] <= 32'd6514;
		word[15'd7439] <= 32'd6515;
		word[15'd7440] <= 32'd6516;
		word[15'd7441] <= 32'd6517;
		word[15'd7442] <= 32'd6518;
		word[15'd7443] <= 32'd6519;
		word[15'd7444] <= 32'd6520;
		word[15'd7445] <= 32'd6521;
		word[15'd7446] <= 32'd6522;
		word[15'd7447] <= 32'd6523;
		word[15'd7448] <= 32'd6524;
		word[15'd7449] <= 32'd6525;
		word[15'd7450] <= 32'd6526;
		word[15'd7451] <= 32'd6527;
		word[15'd7452] <= 32'd6528;
		word[15'd7453] <= 32'd6529;
		word[15'd7454] <= 32'd6530;
		word[15'd7455] <= 32'd6531;
		word[15'd7456] <= 32'd6532;
		word[15'd7457] <= 32'd6533;
		word[15'd7458] <= 32'd6534;
		word[15'd7459] <= 32'd6535;
		word[15'd7460] <= 32'd6536;
		word[15'd7461] <= 32'd6537;
		word[15'd7462] <= 32'd6538;
		word[15'd7463] <= 32'd6539;
		word[15'd7464] <= 32'd6540;
		word[15'd7465] <= 32'd6541;
		word[15'd7466] <= 32'd6542;
		word[15'd7467] <= 32'd6543;
		word[15'd7468] <= 32'd6544;
		word[15'd7469] <= 32'd6545;
		word[15'd7470] <= 32'd6546;
		word[15'd7471] <= 32'd6547;
		word[15'd7472] <= 32'd6548;
		word[15'd7473] <= 32'd6549;
		word[15'd7474] <= 32'd6550;
		word[15'd7475] <= 32'd6551;
		word[15'd7476] <= 32'd6552;
		word[15'd7477] <= 32'd6553;
		word[15'd7478] <= 32'd6554;
		word[15'd7479] <= 32'd6555;
		word[15'd7480] <= 32'd6556;
		word[15'd7481] <= 32'd6557;
		word[15'd7482] <= 32'd6558;
		word[15'd7483] <= 32'd6559;
		word[15'd7484] <= 32'd6560;
		word[15'd7485] <= 32'd6561;
		word[15'd7486] <= 32'd6562;
		word[15'd7487] <= 32'd6563;
		word[15'd7488] <= 32'd6564;
		word[15'd7489] <= 32'd6565;
		word[15'd7490] <= 32'd6566;
		word[15'd7491] <= 32'd6567;
		word[15'd7492] <= 32'd6568;
		word[15'd7493] <= 32'd6569;
		word[15'd7494] <= 32'd6570;
		word[15'd7495] <= 32'd6571;
		word[15'd7496] <= 32'd6572;
		word[15'd7497] <= 32'd6573;
		word[15'd7498] <= 32'd6574;
		word[15'd7499] <= 32'd6575;
		word[15'd7500] <= 32'd6576;
		word[15'd7501] <= 32'd6577;
		word[15'd7502] <= 32'd6578;
		word[15'd7503] <= 32'd6579;
		word[15'd7504] <= 32'd6580;
		word[15'd7505] <= 32'd6581;
		word[15'd7506] <= 32'd6582;
		word[15'd7507] <= 32'd6583;
		word[15'd7508] <= 32'd6584;
		word[15'd7509] <= 32'd6585;
		word[15'd7510] <= 32'd6586;
		word[15'd7511] <= 32'd6587;
		word[15'd7512] <= 32'd6588;
		word[15'd7513] <= 32'd6589;
		word[15'd7514] <= 32'd6590;
		word[15'd7515] <= 32'd6591;
		word[15'd7516] <= 32'd6592;
		word[15'd7517] <= 32'd6593;
		word[15'd7518] <= 32'd6594;
		word[15'd7519] <= 32'd6595;
		word[15'd7520] <= 32'd6596;
		word[15'd7521] <= 32'd6597;
		word[15'd7522] <= 32'd6598;
		word[15'd7523] <= 32'd6599;
		word[15'd7524] <= 32'd6600;
		word[15'd7525] <= 32'd6601;
		word[15'd7526] <= 32'd6602;
		word[15'd7527] <= 32'd6603;
		word[15'd7528] <= 32'd6604;
		word[15'd7529] <= 32'd6605;
		word[15'd7530] <= 32'd6606;
		word[15'd7531] <= 32'd6607;
		word[15'd7532] <= 32'd6608;
		word[15'd7533] <= 32'd6609;
		word[15'd7534] <= 32'd6610;
		word[15'd7535] <= 32'd6611;
		word[15'd7536] <= 32'd6612;
		word[15'd7537] <= 32'd6613;
		word[15'd7538] <= 32'd6614;
		word[15'd7539] <= 32'd6615;
		word[15'd7540] <= 32'd6616;
		word[15'd7541] <= 32'd6617;
		word[15'd7542] <= 32'd6618;
		word[15'd7543] <= 32'd6619;
		word[15'd7544] <= 32'd6620;
		word[15'd7545] <= 32'd6621;
		word[15'd7546] <= 32'd6622;
		word[15'd7547] <= 32'd6623;
		word[15'd7548] <= 32'd6624;
		word[15'd7549] <= 32'd6625;
		word[15'd7550] <= 32'd6626;
		word[15'd7551] <= 32'd6627;
		word[15'd7552] <= 32'd6628;
		word[15'd7553] <= 32'd6629;
		word[15'd7554] <= 32'd6630;
		word[15'd7555] <= 32'd6631;
		word[15'd7556] <= 32'd6632;
		word[15'd7557] <= 32'd6633;
		word[15'd7558] <= 32'd6634;
		word[15'd7559] <= 32'd6635;
		word[15'd7560] <= 32'd6636;
		word[15'd7561] <= 32'd6637;
		word[15'd7562] <= 32'd6638;
		word[15'd7563] <= 32'd6639;
		word[15'd7564] <= 32'd6640;
		word[15'd7565] <= 32'd6641;
		word[15'd7566] <= 32'd6642;
		word[15'd7567] <= 32'd6643;
		word[15'd7568] <= 32'd6644;
		word[15'd7569] <= 32'd6645;
		word[15'd7570] <= 32'd6646;
		word[15'd7571] <= 32'd6647;
		word[15'd7572] <= 32'd6648;
		word[15'd7573] <= 32'd6649;
		word[15'd7574] <= 32'd6650;
		word[15'd7575] <= 32'd6651;
		word[15'd7576] <= 32'd6652;
		word[15'd7577] <= 32'd6653;
		word[15'd7578] <= 32'd6654;
		word[15'd7579] <= 32'd6655;
		word[15'd7580] <= 32'd6656;
		word[15'd7581] <= 32'd6657;
		word[15'd7582] <= 32'd6658;
		word[15'd7583] <= 32'd6659;
		word[15'd7584] <= 32'd6660;
		word[15'd7585] <= 32'd6661;
		word[15'd7586] <= 32'd6662;
		word[15'd7587] <= 32'd6663;
		word[15'd7588] <= 32'd6664;
		word[15'd7589] <= 32'd6665;
		word[15'd7590] <= 32'd6666;
		word[15'd7591] <= 32'd6667;
		word[15'd7592] <= 32'd6668;
		word[15'd7593] <= 32'd6669;
		word[15'd7594] <= 32'd6670;
		word[15'd7595] <= 32'd6671;
		word[15'd7596] <= 32'd6672;
		word[15'd7597] <= 32'd6673;
		word[15'd7598] <= 32'd6674;
		word[15'd7599] <= 32'd6675;
		word[15'd7600] <= 32'd6676;
		word[15'd7601] <= 32'd6677;
		word[15'd7602] <= 32'd6678;
		word[15'd7603] <= 32'd6679;
		word[15'd7604] <= 32'd6680;
		word[15'd7605] <= 32'd6681;
		word[15'd7606] <= 32'd6682;
		word[15'd7607] <= 32'd6683;
		word[15'd7608] <= 32'd6684;
		word[15'd7609] <= 32'd6685;
		word[15'd7610] <= 32'd6686;
		word[15'd7611] <= 32'd6687;
		word[15'd7612] <= 32'd6688;
		word[15'd7613] <= 32'd6689;
		word[15'd7614] <= 32'd6690;
		word[15'd7615] <= 32'd6691;
		word[15'd7616] <= 32'd6692;
		word[15'd7617] <= 32'd6693;
		word[15'd7618] <= 32'd6694;
		word[15'd7619] <= 32'd6695;
		word[15'd7620] <= 32'd6696;
		word[15'd7621] <= 32'd6697;
		word[15'd7622] <= 32'd6698;
		word[15'd7623] <= 32'd6699;
		word[15'd7624] <= 32'd6700;
		word[15'd7625] <= 32'd6701;
		word[15'd7626] <= 32'd6702;
		word[15'd7627] <= 32'd6703;
		word[15'd7628] <= 32'd6704;
		word[15'd7629] <= 32'd6705;
		word[15'd7630] <= 32'd6706;
		word[15'd7631] <= 32'd6707;
		word[15'd7632] <= 32'd6708;
		word[15'd7633] <= 32'd6709;
		word[15'd7634] <= 32'd6710;
		word[15'd7635] <= 32'd6711;
		word[15'd7636] <= 32'd6712;
		word[15'd7637] <= 32'd6713;
		word[15'd7638] <= 32'd6714;
		word[15'd7639] <= 32'd6715;
		word[15'd7640] <= 32'd6716;
		word[15'd7641] <= 32'd6717;
		word[15'd7642] <= 32'd6718;
		word[15'd7643] <= 32'd6719;
		word[15'd7644] <= 32'd6720;
		word[15'd7645] <= 32'd6721;
		word[15'd7646] <= 32'd6722;
		word[15'd7647] <= 32'd6723;
		word[15'd7648] <= 32'd6724;
		word[15'd7649] <= 32'd6725;
		word[15'd7650] <= 32'd6726;
		word[15'd7651] <= 32'd6727;
		word[15'd7652] <= 32'd6728;
		word[15'd7653] <= 32'd6729;
		word[15'd7654] <= 32'd6730;
		word[15'd7655] <= 32'd6731;
		word[15'd7656] <= 32'd6732;
		word[15'd7657] <= 32'd6733;
		word[15'd7658] <= 32'd6734;
		word[15'd7659] <= 32'd6735;
		word[15'd7660] <= 32'd6736;
		word[15'd7661] <= 32'd6737;
		word[15'd7662] <= 32'd6738;
		word[15'd7663] <= 32'd6739;
		word[15'd7664] <= 32'd6740;
		word[15'd7665] <= 32'd6741;
		word[15'd7666] <= 32'd6742;
		word[15'd7667] <= 32'd6743;
		word[15'd7668] <= 32'd6744;
		word[15'd7669] <= 32'd6745;
		word[15'd7670] <= 32'd6746;
		word[15'd7671] <= 32'd6747;
		word[15'd7672] <= 32'd6748;
		word[15'd7673] <= 32'd6749;
		word[15'd7674] <= 32'd6750;
		word[15'd7675] <= 32'd6751;
		word[15'd7676] <= 32'd6752;
		word[15'd7677] <= 32'd6753;
		word[15'd7678] <= 32'd6754;
		word[15'd7679] <= 32'd6755;
		word[15'd7680] <= 32'd6756;
		word[15'd7681] <= 32'd6757;
		word[15'd7682] <= 32'd6758;
		word[15'd7683] <= 32'd6759;
		word[15'd7684] <= 32'd6760;
		word[15'd7685] <= 32'd6761;
		word[15'd7686] <= 32'd6762;
		word[15'd7687] <= 32'd6763;
		word[15'd7688] <= 32'd6764;
		word[15'd7689] <= 32'd6765;
		word[15'd7690] <= 32'd6766;
		word[15'd7691] <= 32'd6767;
		word[15'd7692] <= 32'd6768;
		word[15'd7693] <= 32'd6769;
		word[15'd7694] <= 32'd6770;
		word[15'd7695] <= 32'd6771;
		word[15'd7696] <= 32'd6772;
		word[15'd7697] <= 32'd6773;
		word[15'd7698] <= 32'd6774;
		word[15'd7699] <= 32'd6775;
		word[15'd7700] <= 32'd6776;
		word[15'd7701] <= 32'd6777;
		word[15'd7702] <= 32'd6778;
		word[15'd7703] <= 32'd6779;
		word[15'd7704] <= 32'd6780;
		word[15'd7705] <= 32'd6781;
		word[15'd7706] <= 32'd6782;
		word[15'd7707] <= 32'd6783;
		word[15'd7708] <= 32'd6784;
		word[15'd7709] <= 32'd6785;
		word[15'd7710] <= 32'd6786;
		word[15'd7711] <= 32'd6787;
		word[15'd7712] <= 32'd6788;
		word[15'd7713] <= 32'd6789;
		word[15'd7714] <= 32'd6790;
		word[15'd7715] <= 32'd6791;
		word[15'd7716] <= 32'd6792;
		word[15'd7717] <= 32'd6793;
		word[15'd7718] <= 32'd6794;
		word[15'd7719] <= 32'd6795;
		word[15'd7720] <= 32'd6796;
		word[15'd7721] <= 32'd6797;
		word[15'd7722] <= 32'd6798;
		word[15'd7723] <= 32'd6799;
		word[15'd7724] <= 32'd6800;
		word[15'd7725] <= 32'd6801;
		word[15'd7726] <= 32'd6802;
		word[15'd7727] <= 32'd6803;
		word[15'd7728] <= 32'd6804;
		word[15'd7729] <= 32'd6805;
		word[15'd7730] <= 32'd6806;
		word[15'd7731] <= 32'd6807;
		word[15'd7732] <= 32'd6808;
		word[15'd7733] <= 32'd6809;
		word[15'd7734] <= 32'd6810;
		word[15'd7735] <= 32'd6811;
		word[15'd7736] <= 32'd6812;
		word[15'd7737] <= 32'd6813;
		word[15'd7738] <= 32'd6814;
		word[15'd7739] <= 32'd6815;
		word[15'd7740] <= 32'd6816;
		word[15'd7741] <= 32'd6817;
		word[15'd7742] <= 32'd6818;
		word[15'd7743] <= 32'd6819;
		word[15'd7744] <= 32'd6820;
		word[15'd7745] <= 32'd6821;
		word[15'd7746] <= 32'd6822;
		word[15'd7747] <= 32'd6823;
		word[15'd7748] <= 32'd6824;
		word[15'd7749] <= 32'd6825;
		word[15'd7750] <= 32'd6826;
		word[15'd7751] <= 32'd6827;
		word[15'd7752] <= 32'd6828;
		word[15'd7753] <= 32'd6829;
		word[15'd7754] <= 32'd6830;
		word[15'd7755] <= 32'd6831;
		word[15'd7756] <= 32'd6832;
		word[15'd7757] <= 32'd6833;
		word[15'd7758] <= 32'd6834;
		word[15'd7759] <= 32'd6835;
		word[15'd7760] <= 32'd6836;
		word[15'd7761] <= 32'd6837;
		word[15'd7762] <= 32'd6838;
		word[15'd7763] <= 32'd6839;
		word[15'd7764] <= 32'd6840;
		word[15'd7765] <= 32'd6841;
		word[15'd7766] <= 32'd6842;
		word[15'd7767] <= 32'd6843;
		word[15'd7768] <= 32'd6844;
		word[15'd7769] <= 32'd6845;
		word[15'd7770] <= 32'd6846;
		word[15'd7771] <= 32'd6847;
		word[15'd7772] <= 32'd6848;
		word[15'd7773] <= 32'd6849;
		word[15'd7774] <= 32'd6850;
		word[15'd7775] <= 32'd6851;
		word[15'd7776] <= 32'd6852;
		word[15'd7777] <= 32'd6853;
		word[15'd7778] <= 32'd6854;
		word[15'd7779] <= 32'd6855;
		word[15'd7780] <= 32'd6856;
		word[15'd7781] <= 32'd6857;
		word[15'd7782] <= 32'd6858;
		word[15'd7783] <= 32'd6859;
		word[15'd7784] <= 32'd6860;
		word[15'd7785] <= 32'd6861;
		word[15'd7786] <= 32'd6862;
		word[15'd7787] <= 32'd6863;
		word[15'd7788] <= 32'd6864;
		word[15'd7789] <= 32'd6865;
		word[15'd7790] <= 32'd6866;
		word[15'd7791] <= 32'd6867;
		word[15'd7792] <= 32'd6868;
		word[15'd7793] <= 32'd6869;
		word[15'd7794] <= 32'd6870;
		word[15'd7795] <= 32'd6871;
		word[15'd7796] <= 32'd6872;
		word[15'd7797] <= 32'd6873;
		word[15'd7798] <= 32'd6874;
		word[15'd7799] <= 32'd6875;
		word[15'd7800] <= 32'd6876;
		word[15'd7801] <= 32'd6877;
		word[15'd7802] <= 32'd6878;
		word[15'd7803] <= 32'd6879;
		word[15'd7804] <= 32'd6880;
		word[15'd7805] <= 32'd6881;
		word[15'd7806] <= 32'd6882;
		word[15'd7807] <= 32'd6883;
		word[15'd7808] <= 32'd6884;
		word[15'd7809] <= 32'd6885;
		word[15'd7810] <= 32'd6886;
		word[15'd7811] <= 32'd6887;
		word[15'd7812] <= 32'd6888;
		word[15'd7813] <= 32'd6889;
		word[15'd7814] <= 32'd6890;
		word[15'd7815] <= 32'd6891;
		word[15'd7816] <= 32'd6892;
		word[15'd7817] <= 32'd6893;
		word[15'd7818] <= 32'd6894;
		word[15'd7819] <= 32'd6895;
		word[15'd7820] <= 32'd6896;
		word[15'd7821] <= 32'd6897;
		word[15'd7822] <= 32'd6898;
		word[15'd7823] <= 32'd6899;
		word[15'd7824] <= 32'd6900;
		word[15'd7825] <= 32'd6901;
		word[15'd7826] <= 32'd6902;
		word[15'd7827] <= 32'd6903;
		word[15'd7828] <= 32'd6904;
		word[15'd7829] <= 32'd6905;
		word[15'd7830] <= 32'd6906;
		word[15'd7831] <= 32'd6907;
		word[15'd7832] <= 32'd6908;
		word[15'd7833] <= 32'd6909;
		word[15'd7834] <= 32'd6910;
		word[15'd7835] <= 32'd6911;
		word[15'd7836] <= 32'd6912;
		word[15'd7837] <= 32'd6913;
		word[15'd7838] <= 32'd6914;
		word[15'd7839] <= 32'd6915;
		word[15'd7840] <= 32'd6916;
		word[15'd7841] <= 32'd6917;
		word[15'd7842] <= 32'd6918;
		word[15'd7843] <= 32'd6919;
		word[15'd7844] <= 32'd6920;
		word[15'd7845] <= 32'd6921;
		word[15'd7846] <= 32'd6922;
		word[15'd7847] <= 32'd6923;
		word[15'd7848] <= 32'd6924;
		word[15'd7849] <= 32'd6925;
		word[15'd7850] <= 32'd6926;
		word[15'd7851] <= 32'd6927;
		word[15'd7852] <= 32'd6928;
		word[15'd7853] <= 32'd6929;
		word[15'd7854] <= 32'd6930;
		word[15'd7855] <= 32'd6931;
		word[15'd7856] <= 32'd6932;
		word[15'd7857] <= 32'd6933;
		word[15'd7858] <= 32'd6934;
		word[15'd7859] <= 32'd6935;
		word[15'd7860] <= 32'd6936;
		word[15'd7861] <= 32'd6937;
		word[15'd7862] <= 32'd6938;
		word[15'd7863] <= 32'd6939;
		word[15'd7864] <= 32'd6940;
		word[15'd7865] <= 32'd6941;
		word[15'd7866] <= 32'd6942;
		word[15'd7867] <= 32'd6943;
		word[15'd7868] <= 32'd6944;
		word[15'd7869] <= 32'd6945;
		word[15'd7870] <= 32'd6946;
		word[15'd7871] <= 32'd6947;
		word[15'd7872] <= 32'd6948;
		word[15'd7873] <= 32'd6949;
		word[15'd7874] <= 32'd6950;
		word[15'd7875] <= 32'd6951;
		word[15'd7876] <= 32'd6952;
		word[15'd7877] <= 32'd6953;
		word[15'd7878] <= 32'd6954;
		word[15'd7879] <= 32'd6955;
		word[15'd7880] <= 32'd6956;
		word[15'd7881] <= 32'd6957;
		word[15'd7882] <= 32'd6958;
		word[15'd7883] <= 32'd6959;
		word[15'd7884] <= 32'd6960;
		word[15'd7885] <= 32'd6961;
		word[15'd7886] <= 32'd6962;
		word[15'd7887] <= 32'd6963;
		word[15'd7888] <= 32'd6964;
		word[15'd7889] <= 32'd6965;
		word[15'd7890] <= 32'd6966;
		word[15'd7891] <= 32'd6967;
		word[15'd7892] <= 32'd6968;
		word[15'd7893] <= 32'd6969;
		word[15'd7894] <= 32'd6970;
		word[15'd7895] <= 32'd6971;
		word[15'd7896] <= 32'd6972;
		word[15'd7897] <= 32'd6973;
		word[15'd7898] <= 32'd6974;
		word[15'd7899] <= 32'd6975;
		word[15'd7900] <= 32'd6976;
		word[15'd7901] <= 32'd6977;
		word[15'd7902] <= 32'd6978;
		word[15'd7903] <= 32'd6979;
		word[15'd7904] <= 32'd6980;
		word[15'd7905] <= 32'd6981;
		word[15'd7906] <= 32'd6982;
		word[15'd7907] <= 32'd6983;
		word[15'd7908] <= 32'd6984;
		word[15'd7909] <= 32'd6985;
		word[15'd7910] <= 32'd6986;
		word[15'd7911] <= 32'd6987;
		word[15'd7912] <= 32'd6988;
		word[15'd7913] <= 32'd6989;
		word[15'd7914] <= 32'd6990;
		word[15'd7915] <= 32'd6991;
		word[15'd7916] <= 32'd6992;
		word[15'd7917] <= 32'd6993;
		word[15'd7918] <= 32'd6994;
		word[15'd7919] <= 32'd6995;
		word[15'd7920] <= 32'd6996;
		word[15'd7921] <= 32'd6997;
		word[15'd7922] <= 32'd6998;
		word[15'd7923] <= 32'd6999;
		word[15'd7924] <= 32'd7000;
		word[15'd7925] <= 32'd7001;
		word[15'd7926] <= 32'd7002;
		word[15'd7927] <= 32'd7003;
		word[15'd7928] <= 32'd7004;
		word[15'd7929] <= 32'd7005;
		word[15'd7930] <= 32'd7006;
		word[15'd7931] <= 32'd7007;
		word[15'd7932] <= 32'd7008;
		word[15'd7933] <= 32'd7009;
		word[15'd7934] <= 32'd7010;
		word[15'd7935] <= 32'd7011;
		word[15'd7936] <= 32'd7012;
		word[15'd7937] <= 32'd7013;
		word[15'd7938] <= 32'd7014;
		word[15'd7939] <= 32'd7015;
		word[15'd7940] <= 32'd7016;
		word[15'd7941] <= 32'd7017;
		word[15'd7942] <= 32'd7018;
		word[15'd7943] <= 32'd7019;
		word[15'd7944] <= 32'd7020;
		word[15'd7945] <= 32'd7021;
		word[15'd7946] <= 32'd7022;
		word[15'd7947] <= 32'd7023;
		word[15'd7948] <= 32'd7024;
		word[15'd7949] <= 32'd7025;
		word[15'd7950] <= 32'd7026;
		word[15'd7951] <= 32'd7027;
		word[15'd7952] <= 32'd7028;
		word[15'd7953] <= 32'd7029;
		word[15'd7954] <= 32'd7030;
		word[15'd7955] <= 32'd7031;
		word[15'd7956] <= 32'd7032;
		word[15'd7957] <= 32'd7033;
		word[15'd7958] <= 32'd7034;
		word[15'd7959] <= 32'd7035;
		word[15'd7960] <= 32'd7036;
		word[15'd7961] <= 32'd7037;
		word[15'd7962] <= 32'd7038;
		word[15'd7963] <= 32'd7039;
		word[15'd7964] <= 32'd7040;
		word[15'd7965] <= 32'd7041;
		word[15'd7966] <= 32'd7042;
		word[15'd7967] <= 32'd7043;
		word[15'd7968] <= 32'd7044;
		word[15'd7969] <= 32'd7045;
		word[15'd7970] <= 32'd7046;
		word[15'd7971] <= 32'd7047;
		word[15'd7972] <= 32'd7048;
		word[15'd7973] <= 32'd7049;
		word[15'd7974] <= 32'd7050;
		word[15'd7975] <= 32'd7051;
		word[15'd7976] <= 32'd7052;
		word[15'd7977] <= 32'd7053;
		word[15'd7978] <= 32'd7054;
		word[15'd7979] <= 32'd7055;
		word[15'd7980] <= 32'd7056;
		word[15'd7981] <= 32'd7057;
		word[15'd7982] <= 32'd7058;
		word[15'd7983] <= 32'd7059;
		word[15'd7984] <= 32'd7060;
		word[15'd7985] <= 32'd7061;
		word[15'd7986] <= 32'd7062;
		word[15'd7987] <= 32'd7063;
		word[15'd7988] <= 32'd7064;
		word[15'd7989] <= 32'd7065;
		word[15'd7990] <= 32'd7066;
		word[15'd7991] <= 32'd7067;
		word[15'd7992] <= 32'd7068;
		word[15'd7993] <= 32'd7069;
		word[15'd7994] <= 32'd7070;
		word[15'd7995] <= 32'd7071;
		word[15'd7996] <= 32'd7072;
		word[15'd7997] <= 32'd7073;
		word[15'd7998] <= 32'd7074;
		word[15'd7999] <= 32'd7075;
		word[15'd8000] <= 32'd7076;
		word[15'd8001] <= 32'd7077;
		word[15'd8002] <= 32'd7078;
		word[15'd8003] <= 32'd7079;
		word[15'd8004] <= 32'd7080;
		word[15'd8005] <= 32'd7081;
		word[15'd8006] <= 32'd7082;
		word[15'd8007] <= 32'd7083;
		word[15'd8008] <= 32'd7084;
		word[15'd8009] <= 32'd7085;
		word[15'd8010] <= 32'd7086;
		word[15'd8011] <= 32'd7087;
		word[15'd8012] <= 32'd7088;
		word[15'd8013] <= 32'd7089;
		word[15'd8014] <= 32'd7090;
		word[15'd8015] <= 32'd7091;
		word[15'd8016] <= 32'd7092;
		word[15'd8017] <= 32'd7093;
		word[15'd8018] <= 32'd7094;
		word[15'd8019] <= 32'd7095;
		word[15'd8020] <= 32'd7096;
		word[15'd8021] <= 32'd7097;
		word[15'd8022] <= 32'd7098;
		word[15'd8023] <= 32'd7099;
		word[15'd8024] <= 32'd7100;
		word[15'd8025] <= 32'd7101;
		word[15'd8026] <= 32'd7102;
		word[15'd8027] <= 32'd7103;
		word[15'd8028] <= 32'd7104;
		word[15'd8029] <= 32'd7105;
		word[15'd8030] <= 32'd7106;
		word[15'd8031] <= 32'd7107;
		word[15'd8032] <= 32'd7108;
		word[15'd8033] <= 32'd7109;
		word[15'd8034] <= 32'd7110;
		word[15'd8035] <= 32'd7111;
		word[15'd8036] <= 32'd7112;
		word[15'd8037] <= 32'd7113;
		word[15'd8038] <= 32'd7114;
		word[15'd8039] <= 32'd7115;
		word[15'd8040] <= 32'd7116;
		word[15'd8041] <= 32'd7117;
		word[15'd8042] <= 32'd7118;
		word[15'd8043] <= 32'd7119;
		word[15'd8044] <= 32'd7120;
		word[15'd8045] <= 32'd7121;
		word[15'd8046] <= 32'd7122;
		word[15'd8047] <= 32'd7123;
		word[15'd8048] <= 32'd7124;
		word[15'd8049] <= 32'd7125;
		word[15'd8050] <= 32'd7126;
		word[15'd8051] <= 32'd7127;
		word[15'd8052] <= 32'd7128;
		word[15'd8053] <= 32'd7129;
		word[15'd8054] <= 32'd7130;
		word[15'd8055] <= 32'd7131;
		word[15'd8056] <= 32'd7132;
		word[15'd8057] <= 32'd7133;
		word[15'd8058] <= 32'd7134;
		word[15'd8059] <= 32'd7135;
		word[15'd8060] <= 32'd7136;
		word[15'd8061] <= 32'd7137;
		word[15'd8062] <= 32'd7138;
		word[15'd8063] <= 32'd7139;
		word[15'd8064] <= 32'd7140;
		word[15'd8065] <= 32'd7141;
		word[15'd8066] <= 32'd7142;
		word[15'd8067] <= 32'd7143;
		word[15'd8068] <= 32'd7144;
		word[15'd8069] <= 32'd7145;
		word[15'd8070] <= 32'd7146;
		word[15'd8071] <= 32'd7147;
		word[15'd8072] <= 32'd7148;
		word[15'd8073] <= 32'd7149;
		word[15'd8074] <= 32'd7150;
		word[15'd8075] <= 32'd7151;
		word[15'd8076] <= 32'd7152;
		word[15'd8077] <= 32'd7153;
		word[15'd8078] <= 32'd7154;
		word[15'd8079] <= 32'd7155;
		word[15'd8080] <= 32'd7156;
		word[15'd8081] <= 32'd7157;
		word[15'd8082] <= 32'd7158;
		word[15'd8083] <= 32'd7159;
		word[15'd8084] <= 32'd7160;
		word[15'd8085] <= 32'd7161;
		word[15'd8086] <= 32'd7162;
		word[15'd8087] <= 32'd7163;
		word[15'd8088] <= 32'd7164;
		word[15'd8089] <= 32'd7165;
		word[15'd8090] <= 32'd7166;
		word[15'd8091] <= 32'd7167;
		word[15'd8092] <= 32'd7168;
		word[15'd8093] <= 32'd7169;
		word[15'd8094] <= 32'd7170;
		word[15'd8095] <= 32'd7171;
		word[15'd8096] <= 32'd7172;
		word[15'd8097] <= 32'd7173;
		word[15'd8098] <= 32'd7174;
		word[15'd8099] <= 32'd7175;
		word[15'd8100] <= 32'd7176;
		word[15'd8101] <= 32'd7177;
		word[15'd8102] <= 32'd7178;
		word[15'd8103] <= 32'd7179;
		word[15'd8104] <= 32'd7180;
		word[15'd8105] <= 32'd7181;
		word[15'd8106] <= 32'd7182;
		word[15'd8107] <= 32'd7183;
		word[15'd8108] <= 32'd7184;
		word[15'd8109] <= 32'd7185;
		word[15'd8110] <= 32'd7186;
		word[15'd8111] <= 32'd7187;
		word[15'd8112] <= 32'd7188;
		word[15'd8113] <= 32'd7189;
		word[15'd8114] <= 32'd7190;
		word[15'd8115] <= 32'd7191;
		word[15'd8116] <= 32'd7192;
		word[15'd8117] <= 32'd7193;
		word[15'd8118] <= 32'd7194;
		word[15'd8119] <= 32'd7195;
		word[15'd8120] <= 32'd7196;
		word[15'd8121] <= 32'd7197;
		word[15'd8122] <= 32'd7198;
		word[15'd8123] <= 32'd7199;
		word[15'd8124] <= 32'd7200;
		word[15'd8125] <= 32'd7201;
		word[15'd8126] <= 32'd7202;
		word[15'd8127] <= 32'd7203;
		word[15'd8128] <= 32'd7204;
		word[15'd8129] <= 32'd7205;
		word[15'd8130] <= 32'd7206;
		word[15'd8131] <= 32'd7207;
		word[15'd8132] <= 32'd7208;
		word[15'd8133] <= 32'd7209;
		word[15'd8134] <= 32'd7210;
		word[15'd8135] <= 32'd7211;
		word[15'd8136] <= 32'd7212;
		word[15'd8137] <= 32'd7213;
		word[15'd8138] <= 32'd7214;
		word[15'd8139] <= 32'd7215;
		word[15'd8140] <= 32'd7216;
		word[15'd8141] <= 32'd7217;
		word[15'd8142] <= 32'd7218;
		word[15'd8143] <= 32'd7219;
		word[15'd8144] <= 32'd7220;
		word[15'd8145] <= 32'd7221;
		word[15'd8146] <= 32'd7222;
		word[15'd8147] <= 32'd7223;
		word[15'd8148] <= 32'd7224;
		word[15'd8149] <= 32'd7225;
		word[15'd8150] <= 32'd7226;
		word[15'd8151] <= 32'd7227;
		word[15'd8152] <= 32'd7228;
		word[15'd8153] <= 32'd7229;
		word[15'd8154] <= 32'd7230;
		word[15'd8155] <= 32'd7231;
		word[15'd8156] <= 32'd7232;
		word[15'd8157] <= 32'd7233;
		word[15'd8158] <= 32'd7234;
		word[15'd8159] <= 32'd7235;
		word[15'd8160] <= 32'd7236;
		word[15'd8161] <= 32'd7237;
		word[15'd8162] <= 32'd7238;
		word[15'd8163] <= 32'd7239;
		word[15'd8164] <= 32'd7240;
		word[15'd8165] <= 32'd7241;
		word[15'd8166] <= 32'd7242;
		word[15'd8167] <= 32'd7243;
		word[15'd8168] <= 32'd7244;
		word[15'd8169] <= 32'd7245;
		word[15'd8170] <= 32'd7246;
		word[15'd8171] <= 32'd7247;
		word[15'd8172] <= 32'd7248;
		word[15'd8173] <= 32'd7249;
		word[15'd8174] <= 32'd7250;
		word[15'd8175] <= 32'd7251;
		word[15'd8176] <= 32'd7252;
		word[15'd8177] <= 32'd7253;
		word[15'd8178] <= 32'd7254;
		word[15'd8179] <= 32'd7255;
		word[15'd8180] <= 32'd7256;
		word[15'd8181] <= 32'd7257;
		word[15'd8182] <= 32'd7258;
		word[15'd8183] <= 32'd7259;
		word[15'd8184] <= 32'd7260;
		word[15'd8185] <= 32'd7261;
		word[15'd8186] <= 32'd7262;
		word[15'd8187] <= 32'd7263;
		word[15'd8188] <= 32'd7264;
		word[15'd8189] <= 32'd7265;
		word[15'd8190] <= 32'd7266;
		word[15'd8191] <= 32'd7267;
		word[15'd8192] <= 32'd7268;
		word[15'd8193] <= 32'd7269;
		word[15'd8194] <= 32'd7270;
		word[15'd8195] <= 32'd7271;
		word[15'd8196] <= 32'd7272;
		word[15'd8197] <= 32'd7273;
		word[15'd8198] <= 32'd7274;
		word[15'd8199] <= 32'd7275;
		word[15'd8200] <= 32'd7276;
		word[15'd8201] <= 32'd7277;
		word[15'd8202] <= 32'd7278;
		word[15'd8203] <= 32'd7279;
		word[15'd8204] <= 32'd7280;
		word[15'd8205] <= 32'd7281;
		word[15'd8206] <= 32'd7282;
		word[15'd8207] <= 32'd7283;
		word[15'd8208] <= 32'd7284;
		word[15'd8209] <= 32'd7285;
		word[15'd8210] <= 32'd7286;
		word[15'd8211] <= 32'd7287;
		word[15'd8212] <= 32'd7288;
		word[15'd8213] <= 32'd7289;
		word[15'd8214] <= 32'd7290;
		word[15'd8215] <= 32'd7291;
		word[15'd8216] <= 32'd7292;
		word[15'd8217] <= 32'd7293;
		word[15'd8218] <= 32'd7294;
		word[15'd8219] <= 32'd7295;
		word[15'd8220] <= 32'd7296;
		word[15'd8221] <= 32'd7297;
		word[15'd8222] <= 32'd7298;
		word[15'd8223] <= 32'd7299;
		word[15'd8224] <= 32'd7300;
		word[15'd8225] <= 32'd7301;
		word[15'd8226] <= 32'd7302;
		word[15'd8227] <= 32'd7303;
		word[15'd8228] <= 32'd7304;
		word[15'd8229] <= 32'd7305;
		word[15'd8230] <= 32'd7306;
		word[15'd8231] <= 32'd7307;
		word[15'd8232] <= 32'd7308;
		word[15'd8233] <= 32'd7309;
		word[15'd8234] <= 32'd7310;
		word[15'd8235] <= 32'd7311;
		word[15'd8236] <= 32'd7312;
		word[15'd8237] <= 32'd7313;
		word[15'd8238] <= 32'd7314;
		word[15'd8239] <= 32'd7315;
		word[15'd8240] <= 32'd7316;
		word[15'd8241] <= 32'd7317;
		word[15'd8242] <= 32'd7318;
		word[15'd8243] <= 32'd7319;
		word[15'd8244] <= 32'd7320;
		word[15'd8245] <= 32'd7321;
		word[15'd8246] <= 32'd7322;
		word[15'd8247] <= 32'd7323;
		word[15'd8248] <= 32'd7324;
		word[15'd8249] <= 32'd7325;
		word[15'd8250] <= 32'd7326;
		word[15'd8251] <= 32'd7327;
		word[15'd8252] <= 32'd7328;
		word[15'd8253] <= 32'd7329;
		word[15'd8254] <= 32'd7330;
		word[15'd8255] <= 32'd7331;
		word[15'd8256] <= 32'd7332;
		word[15'd8257] <= 32'd7333;
		word[15'd8258] <= 32'd7334;
		word[15'd8259] <= 32'd7335;
		word[15'd8260] <= 32'd7336;
		word[15'd8261] <= 32'd7337;
		word[15'd8262] <= 32'd7338;
		word[15'd8263] <= 32'd7339;
		word[15'd8264] <= 32'd7340;
		word[15'd8265] <= 32'd7341;
		word[15'd8266] <= 32'd7342;
		word[15'd8267] <= 32'd7343;
		word[15'd8268] <= 32'd7344;
		word[15'd8269] <= 32'd7345;
		word[15'd8270] <= 32'd7346;
		word[15'd8271] <= 32'd7347;
		word[15'd8272] <= 32'd7348;
		word[15'd8273] <= 32'd7349;
		word[15'd8274] <= 32'd7350;
		word[15'd8275] <= 32'd7351;
		word[15'd8276] <= 32'd7352;
		word[15'd8277] <= 32'd7353;
		word[15'd8278] <= 32'd7354;
		word[15'd8279] <= 32'd7355;
		word[15'd8280] <= 32'd7356;
		word[15'd8281] <= 32'd7357;
		word[15'd8282] <= 32'd7358;
		word[15'd8283] <= 32'd7359;
		word[15'd8284] <= 32'd7360;
		word[15'd8285] <= 32'd7361;
		word[15'd8286] <= 32'd7362;
		word[15'd8287] <= 32'd7363;
		word[15'd8288] <= 32'd7364;
		word[15'd8289] <= 32'd7365;
		word[15'd8290] <= 32'd7366;
		word[15'd8291] <= 32'd7367;
		word[15'd8292] <= 32'd7368;
		word[15'd8293] <= 32'd7369;
		word[15'd8294] <= 32'd7370;
		word[15'd8295] <= 32'd7371;
		word[15'd8296] <= 32'd7372;
		word[15'd8297] <= 32'd7373;
		word[15'd8298] <= 32'd7374;
		word[15'd8299] <= 32'd7375;
		word[15'd8300] <= 32'd7376;
		word[15'd8301] <= 32'd7377;
		word[15'd8302] <= 32'd7378;
		word[15'd8303] <= 32'd7379;
		word[15'd8304] <= 32'd7380;
		word[15'd8305] <= 32'd7381;
		word[15'd8306] <= 32'd7382;
		word[15'd8307] <= 32'd7383;
		word[15'd8308] <= 32'd7384;
		word[15'd8309] <= 32'd7385;
		word[15'd8310] <= 32'd7386;
		word[15'd8311] <= 32'd7387;
		word[15'd8312] <= 32'd7388;
		word[15'd8313] <= 32'd7389;
		word[15'd8314] <= 32'd7390;
		word[15'd8315] <= 32'd7391;
		word[15'd8316] <= 32'd7392;
		word[15'd8317] <= 32'd7393;
		word[15'd8318] <= 32'd7394;
		word[15'd8319] <= 32'd7395;
		word[15'd8320] <= 32'd7396;
		word[15'd8321] <= 32'd7397;
		word[15'd8322] <= 32'd7398;
		word[15'd8323] <= 32'd7399;
		word[15'd8324] <= 32'd7400;
		word[15'd8325] <= 32'd7401;
		word[15'd8326] <= 32'd7402;
		word[15'd8327] <= 32'd7403;
		word[15'd8328] <= 32'd7404;
		word[15'd8329] <= 32'd7405;
		word[15'd8330] <= 32'd7406;
		word[15'd8331] <= 32'd7407;
		word[15'd8332] <= 32'd7408;
		word[15'd8333] <= 32'd7409;
		word[15'd8334] <= 32'd7410;
		word[15'd8335] <= 32'd7411;
		word[15'd8336] <= 32'd7412;
		word[15'd8337] <= 32'd7413;
		word[15'd8338] <= 32'd7414;
		word[15'd8339] <= 32'd7415;
		word[15'd8340] <= 32'd7416;
		word[15'd8341] <= 32'd7417;
		word[15'd8342] <= 32'd7418;
		word[15'd8343] <= 32'd7419;
		word[15'd8344] <= 32'd7420;
		word[15'd8345] <= 32'd7421;
		word[15'd8346] <= 32'd7422;
		word[15'd8347] <= 32'd7423;
		word[15'd8348] <= 32'd7424;
		word[15'd8349] <= 32'd7425;
		word[15'd8350] <= 32'd7426;
		word[15'd8351] <= 32'd7427;
		word[15'd8352] <= 32'd7428;
		word[15'd8353] <= 32'd7429;
		word[15'd8354] <= 32'd7430;
		word[15'd8355] <= 32'd7431;
		word[15'd8356] <= 32'd7432;
		word[15'd8357] <= 32'd7433;
		word[15'd8358] <= 32'd7434;
		word[15'd8359] <= 32'd7435;
		word[15'd8360] <= 32'd7436;
		word[15'd8361] <= 32'd7437;
		word[15'd8362] <= 32'd7438;
		word[15'd8363] <= 32'd7439;
		word[15'd8364] <= 32'd7440;
		word[15'd8365] <= 32'd7441;
		word[15'd8366] <= 32'd7442;
		word[15'd8367] <= 32'd7443;
		word[15'd8368] <= 32'd7444;
		word[15'd8369] <= 32'd7445;
		word[15'd8370] <= 32'd7446;
		word[15'd8371] <= 32'd7447;
		word[15'd8372] <= 32'd7448;
		word[15'd8373] <= 32'd7449;
		word[15'd8374] <= 32'd7450;
		word[15'd8375] <= 32'd7451;
		word[15'd8376] <= 32'd7452;
		word[15'd8377] <= 32'd7453;
		word[15'd8378] <= 32'd7454;
		word[15'd8379] <= 32'd7455;
		word[15'd8380] <= 32'd7456;
		word[15'd8381] <= 32'd7457;
		word[15'd8382] <= 32'd7458;
		word[15'd8383] <= 32'd7459;
		word[15'd8384] <= 32'd7460;
		word[15'd8385] <= 32'd7461;
		word[15'd8386] <= 32'd7462;
		word[15'd8387] <= 32'd7463;
		word[15'd8388] <= 32'd7464;
		word[15'd8389] <= 32'd7465;
		word[15'd8390] <= 32'd7466;
		word[15'd8391] <= 32'd7467;
		word[15'd8392] <= 32'd7468;
		word[15'd8393] <= 32'd7469;
		word[15'd8394] <= 32'd7470;
		word[15'd8395] <= 32'd7471;
		word[15'd8396] <= 32'd7472;
		word[15'd8397] <= 32'd7473;
		word[15'd8398] <= 32'd7474;
		word[15'd8399] <= 32'd7475;
		word[15'd8400] <= 32'd7476;
		word[15'd8401] <= 32'd7477;
		word[15'd8402] <= 32'd7478;
		word[15'd8403] <= 32'd7479;
		word[15'd8404] <= 32'd7480;
		word[15'd8405] <= 32'd7481;
		word[15'd8406] <= 32'd7482;
		word[15'd8407] <= 32'd7483;
		word[15'd8408] <= 32'd7484;
		word[15'd8409] <= 32'd7485;
		word[15'd8410] <= 32'd7486;
		word[15'd8411] <= 32'd7487;
		word[15'd8412] <= 32'd7488;
		word[15'd8413] <= 32'd7489;
		word[15'd8414] <= 32'd7490;
		word[15'd8415] <= 32'd7491;
		word[15'd8416] <= 32'd7492;
		word[15'd8417] <= 32'd7493;
		word[15'd8418] <= 32'd7494;
		word[15'd8419] <= 32'd7495;
		word[15'd8420] <= 32'd7496;
		word[15'd8421] <= 32'd7497;
		word[15'd8422] <= 32'd7498;
		word[15'd8423] <= 32'd7499;
		word[15'd8424] <= 32'd7500;
		word[15'd8425] <= 32'd7501;
		word[15'd8426] <= 32'd7502;
		word[15'd8427] <= 32'd7503;
		word[15'd8428] <= 32'd7504;
		word[15'd8429] <= 32'd7505;
		word[15'd8430] <= 32'd7506;
		word[15'd8431] <= 32'd7507;
		word[15'd8432] <= 32'd7508;
		word[15'd8433] <= 32'd7509;
		word[15'd8434] <= 32'd7510;
		word[15'd8435] <= 32'd7511;
		word[15'd8436] <= 32'd7512;
		word[15'd8437] <= 32'd7513;
		word[15'd8438] <= 32'd7514;
		word[15'd8439] <= 32'd7515;
		word[15'd8440] <= 32'd7516;
		word[15'd8441] <= 32'd7517;
		word[15'd8442] <= 32'd7518;
		word[15'd8443] <= 32'd7519;
		word[15'd8444] <= 32'd7520;
		word[15'd8445] <= 32'd7521;
		word[15'd8446] <= 32'd7522;
		word[15'd8447] <= 32'd7523;
		word[15'd8448] <= 32'd7524;
		word[15'd8449] <= 32'd7525;
		word[15'd8450] <= 32'd7526;
		word[15'd8451] <= 32'd7527;
		word[15'd8452] <= 32'd7528;
		word[15'd8453] <= 32'd7529;
		word[15'd8454] <= 32'd7530;
		word[15'd8455] <= 32'd7531;
		word[15'd8456] <= 32'd7532;
		word[15'd8457] <= 32'd7533;
		word[15'd8458] <= 32'd7534;
		word[15'd8459] <= 32'd7535;
		word[15'd8460] <= 32'd7536;
		word[15'd8461] <= 32'd7537;
		word[15'd8462] <= 32'd7538;
		word[15'd8463] <= 32'd7539;
		word[15'd8464] <= 32'd7540;
		word[15'd8465] <= 32'd7541;
		word[15'd8466] <= 32'd7542;
		word[15'd8467] <= 32'd7543;
		word[15'd8468] <= 32'd7544;
		word[15'd8469] <= 32'd7545;
		word[15'd8470] <= 32'd7546;
		word[15'd8471] <= 32'd7547;
		word[15'd8472] <= 32'd7548;
		word[15'd8473] <= 32'd7549;
		word[15'd8474] <= 32'd7550;
		word[15'd8475] <= 32'd7551;
		word[15'd8476] <= 32'd7552;
		word[15'd8477] <= 32'd7553;
		word[15'd8478] <= 32'd7554;
		word[15'd8479] <= 32'd7555;
		word[15'd8480] <= 32'd7556;
		word[15'd8481] <= 32'd7557;
		word[15'd8482] <= 32'd7558;
		word[15'd8483] <= 32'd7559;
		word[15'd8484] <= 32'd7560;
		word[15'd8485] <= 32'd7561;
		word[15'd8486] <= 32'd7562;
		word[15'd8487] <= 32'd7563;
		word[15'd8488] <= 32'd7564;
		word[15'd8489] <= 32'd7565;
		word[15'd8490] <= 32'd7566;
		word[15'd8491] <= 32'd7567;
		word[15'd8492] <= 32'd7568;
		word[15'd8493] <= 32'd7569;
		word[15'd8494] <= 32'd7570;
		word[15'd8495] <= 32'd7571;
		word[15'd8496] <= 32'd7572;
		word[15'd8497] <= 32'd7573;
		word[15'd8498] <= 32'd7574;
		word[15'd8499] <= 32'd7575;
		word[15'd8500] <= 32'd7576;
		word[15'd8501] <= 32'd7577;
		word[15'd8502] <= 32'd7578;
		word[15'd8503] <= 32'd7579;
		word[15'd8504] <= 32'd7580;
		word[15'd8505] <= 32'd7581;
		word[15'd8506] <= 32'd7582;
		word[15'd8507] <= 32'd7583;
		word[15'd8508] <= 32'd7584;
		word[15'd8509] <= 32'd7585;
		word[15'd8510] <= 32'd7586;
		word[15'd8511] <= 32'd7587;
		word[15'd8512] <= 32'd7588;
		word[15'd8513] <= 32'd7589;
		word[15'd8514] <= 32'd7590;
		word[15'd8515] <= 32'd7591;
		word[15'd8516] <= 32'd7592;
		word[15'd8517] <= 32'd7593;
		word[15'd8518] <= 32'd7594;
		word[15'd8519] <= 32'd7595;
		word[15'd8520] <= 32'd7596;
		word[15'd8521] <= 32'd7597;
		word[15'd8522] <= 32'd7598;
		word[15'd8523] <= 32'd7599;
		word[15'd8524] <= 32'd7600;
		word[15'd8525] <= 32'd7601;
		word[15'd8526] <= 32'd7602;
		word[15'd8527] <= 32'd7603;
		word[15'd8528] <= 32'd7604;
		word[15'd8529] <= 32'd7605;
		word[15'd8530] <= 32'd7606;
		word[15'd8531] <= 32'd7607;
		word[15'd8532] <= 32'd7608;
		word[15'd8533] <= 32'd7609;
		word[15'd8534] <= 32'd7610;
		word[15'd8535] <= 32'd7611;
		word[15'd8536] <= 32'd7612;
		word[15'd8537] <= 32'd7613;
		word[15'd8538] <= 32'd7614;
		word[15'd8539] <= 32'd7615;
		word[15'd8540] <= 32'd7616;
		word[15'd8541] <= 32'd7617;
		word[15'd8542] <= 32'd7618;
		word[15'd8543] <= 32'd7619;
		word[15'd8544] <= 32'd7620;
		word[15'd8545] <= 32'd7621;
		word[15'd8546] <= 32'd7622;
		word[15'd8547] <= 32'd7623;
		word[15'd8548] <= 32'd7624;
		word[15'd8549] <= 32'd7625;
		word[15'd8550] <= 32'd7626;
		word[15'd8551] <= 32'd7627;
		word[15'd8552] <= 32'd7628;
		word[15'd8553] <= 32'd7629;
		word[15'd8554] <= 32'd7630;
		word[15'd8555] <= 32'd7631;
		word[15'd8556] <= 32'd7632;
		word[15'd8557] <= 32'd7633;
		word[15'd8558] <= 32'd7634;
		word[15'd8559] <= 32'd7635;
		word[15'd8560] <= 32'd7636;
		word[15'd8561] <= 32'd7637;
		word[15'd8562] <= 32'd7638;
		word[15'd8563] <= 32'd7639;
		word[15'd8564] <= 32'd7640;
		word[15'd8565] <= 32'd7641;
		word[15'd8566] <= 32'd7642;
		word[15'd8567] <= 32'd7643;
		word[15'd8568] <= 32'd7644;
		word[15'd8569] <= 32'd7645;
		word[15'd8570] <= 32'd7646;
		word[15'd8571] <= 32'd7647;
		word[15'd8572] <= 32'd7648;
		word[15'd8573] <= 32'd7649;
		word[15'd8574] <= 32'd7650;
		word[15'd8575] <= 32'd7651;
		word[15'd8576] <= 32'd7652;
		word[15'd8577] <= 32'd7653;
		word[15'd8578] <= 32'd7654;
		word[15'd8579] <= 32'd7655;
		word[15'd8580] <= 32'd7656;
		word[15'd8581] <= 32'd7657;
		word[15'd8582] <= 32'd7658;
		word[15'd8583] <= 32'd7659;
		word[15'd8584] <= 32'd7660;
		word[15'd8585] <= 32'd7661;
		word[15'd8586] <= 32'd7662;
		word[15'd8587] <= 32'd7663;
		word[15'd8588] <= 32'd7664;
		word[15'd8589] <= 32'd7665;
		word[15'd8590] <= 32'd7666;
		word[15'd8591] <= 32'd7667;
		word[15'd8592] <= 32'd7668;
		word[15'd8593] <= 32'd7669;
		word[15'd8594] <= 32'd7670;
		word[15'd8595] <= 32'd7671;
		word[15'd8596] <= 32'd7672;
		word[15'd8597] <= 32'd7673;
		word[15'd8598] <= 32'd7674;
		word[15'd8599] <= 32'd7675;
		word[15'd8600] <= 32'd7676;
		word[15'd8601] <= 32'd7677;
		word[15'd8602] <= 32'd7678;
		word[15'd8603] <= 32'd7679;
		word[15'd8604] <= 32'd7680;
		word[15'd8605] <= 32'd7681;
		word[15'd8606] <= 32'd7682;
		word[15'd8607] <= 32'd7683;
		word[15'd8608] <= 32'd7684;
		word[15'd8609] <= 32'd7685;
		word[15'd8610] <= 32'd7686;
		word[15'd8611] <= 32'd7687;
		word[15'd8612] <= 32'd7688;
		word[15'd8613] <= 32'd7689;
		word[15'd8614] <= 32'd7690;
		word[15'd8615] <= 32'd7691;
		word[15'd8616] <= 32'd7692;
		word[15'd8617] <= 32'd7693;
		word[15'd8618] <= 32'd7694;
		word[15'd8619] <= 32'd7695;
		word[15'd8620] <= 32'd7696;
		word[15'd8621] <= 32'd7697;
		word[15'd8622] <= 32'd7698;
		word[15'd8623] <= 32'd7699;
		word[15'd8624] <= 32'd7700;
		word[15'd8625] <= 32'd7701;
		word[15'd8626] <= 32'd7702;
		word[15'd8627] <= 32'd7703;
		word[15'd8628] <= 32'd7704;
		word[15'd8629] <= 32'd7705;
		word[15'd8630] <= 32'd7706;
		word[15'd8631] <= 32'd7707;
		word[15'd8632] <= 32'd7708;
		word[15'd8633] <= 32'd7709;
		word[15'd8634] <= 32'd7710;
		word[15'd8635] <= 32'd7711;
		word[15'd8636] <= 32'd7712;
		word[15'd8637] <= 32'd7713;
		word[15'd8638] <= 32'd7714;
		word[15'd8639] <= 32'd7715;
		word[15'd8640] <= 32'd7716;
		word[15'd8641] <= 32'd7717;
		word[15'd8642] <= 32'd7718;
		word[15'd8643] <= 32'd7719;
		word[15'd8644] <= 32'd7720;
		word[15'd8645] <= 32'd7721;
		word[15'd8646] <= 32'd7722;
		word[15'd8647] <= 32'd7723;
		word[15'd8648] <= 32'd7724;
		word[15'd8649] <= 32'd7725;
		word[15'd8650] <= 32'd7726;
		word[15'd8651] <= 32'd7727;
		word[15'd8652] <= 32'd7728;
		word[15'd8653] <= 32'd7729;
		word[15'd8654] <= 32'd7730;
		word[15'd8655] <= 32'd7731;
		word[15'd8656] <= 32'd7732;
		word[15'd8657] <= 32'd7733;
		word[15'd8658] <= 32'd7734;
		word[15'd8659] <= 32'd7735;
		word[15'd8660] <= 32'd7736;
		word[15'd8661] <= 32'd7737;
		word[15'd8662] <= 32'd7738;
		word[15'd8663] <= 32'd7739;
		word[15'd8664] <= 32'd7740;
		word[15'd8665] <= 32'd7741;
		word[15'd8666] <= 32'd7742;
		word[15'd8667] <= 32'd7743;
		word[15'd8668] <= 32'd7744;
		word[15'd8669] <= 32'd7745;
		word[15'd8670] <= 32'd7746;
		word[15'd8671] <= 32'd7747;
		word[15'd8672] <= 32'd7748;
		word[15'd8673] <= 32'd7749;
		word[15'd8674] <= 32'd7750;
		word[15'd8675] <= 32'd7751;
		word[15'd8676] <= 32'd7752;
		word[15'd8677] <= 32'd7753;
		word[15'd8678] <= 32'd7754;
		word[15'd8679] <= 32'd7755;
		word[15'd8680] <= 32'd7756;
		word[15'd8681] <= 32'd7757;
		word[15'd8682] <= 32'd7758;
		word[15'd8683] <= 32'd7759;
		word[15'd8684] <= 32'd7760;
		word[15'd8685] <= 32'd7761;
		word[15'd8686] <= 32'd7762;
		word[15'd8687] <= 32'd7763;
		word[15'd8688] <= 32'd7764;
		word[15'd8689] <= 32'd7765;
		word[15'd8690] <= 32'd7766;
		word[15'd8691] <= 32'd7767;
		word[15'd8692] <= 32'd7768;
		word[15'd8693] <= 32'd7769;
		word[15'd8694] <= 32'd7770;
		word[15'd8695] <= 32'd7771;
		word[15'd8696] <= 32'd7772;
		word[15'd8697] <= 32'd7773;
		word[15'd8698] <= 32'd7774;
		word[15'd8699] <= 32'd7775;
		word[15'd8700] <= 32'd7776;
		word[15'd8701] <= 32'd7777;
		word[15'd8702] <= 32'd7778;
		word[15'd8703] <= 32'd7779;
		word[15'd8704] <= 32'd7780;
		word[15'd8705] <= 32'd7781;
		word[15'd8706] <= 32'd7782;
		word[15'd8707] <= 32'd7783;
		word[15'd8708] <= 32'd7784;
		word[15'd8709] <= 32'd7785;
		word[15'd8710] <= 32'd7786;
		word[15'd8711] <= 32'd7787;
		word[15'd8712] <= 32'd7788;
		word[15'd8713] <= 32'd7789;
		word[15'd8714] <= 32'd7790;
		word[15'd8715] <= 32'd7791;
		word[15'd8716] <= 32'd7792;
		word[15'd8717] <= 32'd7793;
		word[15'd8718] <= 32'd7794;
		word[15'd8719] <= 32'd7795;
		word[15'd8720] <= 32'd7796;
		word[15'd8721] <= 32'd7797;
		word[15'd8722] <= 32'd7798;
		word[15'd8723] <= 32'd7799;
		word[15'd8724] <= 32'd7800;
		word[15'd8725] <= 32'd7801;
		word[15'd8726] <= 32'd7802;
		word[15'd8727] <= 32'd7803;
		word[15'd8728] <= 32'd7804;
		word[15'd8729] <= 32'd7805;
		word[15'd8730] <= 32'd7806;
		word[15'd8731] <= 32'd7807;
		word[15'd8732] <= 32'd7808;
		word[15'd8733] <= 32'd7809;
		word[15'd8734] <= 32'd7810;
		word[15'd8735] <= 32'd7811;
		word[15'd8736] <= 32'd7812;
		word[15'd8737] <= 32'd7813;
		word[15'd8738] <= 32'd7814;
		word[15'd8739] <= 32'd7815;
		word[15'd8740] <= 32'd7816;
		word[15'd8741] <= 32'd7817;
		word[15'd8742] <= 32'd7818;
		word[15'd8743] <= 32'd7819;
		word[15'd8744] <= 32'd7820;
		word[15'd8745] <= 32'd7821;
		word[15'd8746] <= 32'd7822;
		word[15'd8747] <= 32'd7823;
		word[15'd8748] <= 32'd7824;
		word[15'd8749] <= 32'd7825;
		word[15'd8750] <= 32'd7826;
		word[15'd8751] <= 32'd7827;
		word[15'd8752] <= 32'd7828;
		word[15'd8753] <= 32'd7829;
		word[15'd8754] <= 32'd7830;
		word[15'd8755] <= 32'd7831;
		word[15'd8756] <= 32'd7832;
		word[15'd8757] <= 32'd7833;
		word[15'd8758] <= 32'd7834;
		word[15'd8759] <= 32'd7835;
		word[15'd8760] <= 32'd7836;
		word[15'd8761] <= 32'd7837;
		word[15'd8762] <= 32'd7838;
		word[15'd8763] <= 32'd7839;
		word[15'd8764] <= 32'd7840;
		word[15'd8765] <= 32'd7841;
		word[15'd8766] <= 32'd7842;
		word[15'd8767] <= 32'd7843;
		word[15'd8768] <= 32'd7844;
		word[15'd8769] <= 32'd7845;
		word[15'd8770] <= 32'd7846;
		word[15'd8771] <= 32'd7847;
		word[15'd8772] <= 32'd7848;
		word[15'd8773] <= 32'd7849;
		word[15'd8774] <= 32'd7850;
		word[15'd8775] <= 32'd7851;
		word[15'd8776] <= 32'd7852;
		word[15'd8777] <= 32'd7853;
		word[15'd8778] <= 32'd7854;
		word[15'd8779] <= 32'd7855;
		word[15'd8780] <= 32'd7856;
		word[15'd8781] <= 32'd7857;
		word[15'd8782] <= 32'd7858;
		word[15'd8783] <= 32'd7859;
		word[15'd8784] <= 32'd7860;
		word[15'd8785] <= 32'd7861;
		word[15'd8786] <= 32'd7862;
		word[15'd8787] <= 32'd7863;
		word[15'd8788] <= 32'd7864;
		word[15'd8789] <= 32'd7865;
		word[15'd8790] <= 32'd7866;
		word[15'd8791] <= 32'd7867;
		word[15'd8792] <= 32'd7868;
		word[15'd8793] <= 32'd7869;
		word[15'd8794] <= 32'd7870;
		word[15'd8795] <= 32'd7871;
		word[15'd8796] <= 32'd7872;
		word[15'd8797] <= 32'd7873;
		word[15'd8798] <= 32'd7874;
		word[15'd8799] <= 32'd7875;
		word[15'd8800] <= 32'd7876;
		word[15'd8801] <= 32'd7877;
		word[15'd8802] <= 32'd7878;
		word[15'd8803] <= 32'd7879;
		word[15'd8804] <= 32'd7880;
		word[15'd8805] <= 32'd7881;
		word[15'd8806] <= 32'd7882;
		word[15'd8807] <= 32'd7883;
		word[15'd8808] <= 32'd7884;
		word[15'd8809] <= 32'd7885;
		word[15'd8810] <= 32'd7886;
		word[15'd8811] <= 32'd7887;
		word[15'd8812] <= 32'd7888;
		word[15'd8813] <= 32'd7889;
		word[15'd8814] <= 32'd7890;
		word[15'd8815] <= 32'd7891;
		word[15'd8816] <= 32'd7892;
		word[15'd8817] <= 32'd7893;
		word[15'd8818] <= 32'd7894;
		word[15'd8819] <= 32'd7895;
		word[15'd8820] <= 32'd7896;
		word[15'd8821] <= 32'd7897;
		word[15'd8822] <= 32'd7898;
		word[15'd8823] <= 32'd7899;
		word[15'd8824] <= 32'd7900;
		word[15'd8825] <= 32'd7901;
		word[15'd8826] <= 32'd7902;
		word[15'd8827] <= 32'd7903;
		word[15'd8828] <= 32'd7904;
		word[15'd8829] <= 32'd7905;
		word[15'd8830] <= 32'd7906;
		word[15'd8831] <= 32'd7907;
		word[15'd8832] <= 32'd7908;
		word[15'd8833] <= 32'd7909;
		word[15'd8834] <= 32'd7910;
		word[15'd8835] <= 32'd7911;
		word[15'd8836] <= 32'd7912;
		word[15'd8837] <= 32'd7913;
		word[15'd8838] <= 32'd7914;
		word[15'd8839] <= 32'd7915;
		word[15'd8840] <= 32'd7916;
		word[15'd8841] <= 32'd7917;
		word[15'd8842] <= 32'd7918;
		word[15'd8843] <= 32'd7919;
		word[15'd8844] <= 32'd7920;
		word[15'd8845] <= 32'd7921;
		word[15'd8846] <= 32'd7922;
		word[15'd8847] <= 32'd7923;
		word[15'd8848] <= 32'd7924;
		word[15'd8849] <= 32'd7925;
		word[15'd8850] <= 32'd7926;
		word[15'd8851] <= 32'd7927;
		word[15'd8852] <= 32'd7928;
		word[15'd8853] <= 32'd7929;
		word[15'd8854] <= 32'd7930;
		word[15'd8855] <= 32'd7931;
		word[15'd8856] <= 32'd7932;
		word[15'd8857] <= 32'd7933;
		word[15'd8858] <= 32'd7934;
		word[15'd8859] <= 32'd7935;
		word[15'd8860] <= 32'd7936;
		word[15'd8861] <= 32'd7937;
		word[15'd8862] <= 32'd7938;
		word[15'd8863] <= 32'd7939;
		word[15'd8864] <= 32'd7940;
		word[15'd8865] <= 32'd7941;
		word[15'd8866] <= 32'd7942;
		word[15'd8867] <= 32'd7943;
		word[15'd8868] <= 32'd7944;
		word[15'd8869] <= 32'd7945;
		word[15'd8870] <= 32'd7946;
		word[15'd8871] <= 32'd7947;
		word[15'd8872] <= 32'd7948;
		word[15'd8873] <= 32'd7949;
		word[15'd8874] <= 32'd7950;
		word[15'd8875] <= 32'd7951;
		word[15'd8876] <= 32'd7952;
		word[15'd8877] <= 32'd7953;
		word[15'd8878] <= 32'd7954;
		word[15'd8879] <= 32'd7955;
		word[15'd8880] <= 32'd7956;
		word[15'd8881] <= 32'd7957;
		word[15'd8882] <= 32'd7958;
		word[15'd8883] <= 32'd7959;
		word[15'd8884] <= 32'd7960;
		word[15'd8885] <= 32'd7961;
		word[15'd8886] <= 32'd7962;
		word[15'd8887] <= 32'd7963;
		word[15'd8888] <= 32'd7964;
		word[15'd8889] <= 32'd7965;
		word[15'd8890] <= 32'd7966;
		word[15'd8891] <= 32'd7967;
		word[15'd8892] <= 32'd7968;
		word[15'd8893] <= 32'd7969;
		word[15'd8894] <= 32'd7970;
		word[15'd8895] <= 32'd7971;
		word[15'd8896] <= 32'd7972;
		word[15'd8897] <= 32'd7973;
		word[15'd8898] <= 32'd7974;
		word[15'd8899] <= 32'd7975;
		word[15'd8900] <= 32'd7976;
		word[15'd8901] <= 32'd7977;
		word[15'd8902] <= 32'd7978;
		word[15'd8903] <= 32'd7979;
		word[15'd8904] <= 32'd7980;
		word[15'd8905] <= 32'd7981;
		word[15'd8906] <= 32'd7982;
		word[15'd8907] <= 32'd7983;
		word[15'd8908] <= 32'd7984;
		word[15'd8909] <= 32'd7985;
		word[15'd8910] <= 32'd7986;
		word[15'd8911] <= 32'd7987;
		word[15'd8912] <= 32'd7988;
		word[15'd8913] <= 32'd7989;
		word[15'd8914] <= 32'd7990;
		word[15'd8915] <= 32'd7991;
		word[15'd8916] <= 32'd7992;
		word[15'd8917] <= 32'd7993;
		word[15'd8918] <= 32'd7994;
		word[15'd8919] <= 32'd7995;
		word[15'd8920] <= 32'd7996;
		word[15'd8921] <= 32'd7997;
		word[15'd8922] <= 32'd7998;
		word[15'd8923] <= 32'd7999;
		word[15'd8924] <= 32'd8000;
		word[15'd8925] <= 32'd8001;
		word[15'd8926] <= 32'd8002;
		word[15'd8927] <= 32'd8003;
		word[15'd8928] <= 32'd8004;
		word[15'd8929] <= 32'd8005;
		word[15'd8930] <= 32'd8006;
		word[15'd8931] <= 32'd8007;
		word[15'd8932] <= 32'd8008;
		word[15'd8933] <= 32'd8009;
		word[15'd8934] <= 32'd8010;
		word[15'd8935] <= 32'd8011;
		word[15'd8936] <= 32'd8012;
		word[15'd8937] <= 32'd8013;
		word[15'd8938] <= 32'd8014;
		word[15'd8939] <= 32'd8015;
		word[15'd8940] <= 32'd8016;
		word[15'd8941] <= 32'd8017;
		word[15'd8942] <= 32'd8018;
		word[15'd8943] <= 32'd8019;
		word[15'd8944] <= 32'd8020;
		word[15'd8945] <= 32'd8021;
		word[15'd8946] <= 32'd8022;
		word[15'd8947] <= 32'd8023;
		word[15'd8948] <= 32'd8024;
		word[15'd8949] <= 32'd8025;
		word[15'd8950] <= 32'd8026;
		word[15'd8951] <= 32'd8027;
		word[15'd8952] <= 32'd8028;
		word[15'd8953] <= 32'd8029;
		word[15'd8954] <= 32'd8030;
		word[15'd8955] <= 32'd8031;
		word[15'd8956] <= 32'd8032;
		word[15'd8957] <= 32'd8033;
		word[15'd8958] <= 32'd8034;
		word[15'd8959] <= 32'd8035;
		word[15'd8960] <= 32'd8036;
		word[15'd8961] <= 32'd8037;
		word[15'd8962] <= 32'd8038;
		word[15'd8963] <= 32'd8039;
		word[15'd8964] <= 32'd8040;
		word[15'd8965] <= 32'd8041;
		word[15'd8966] <= 32'd8042;
		word[15'd8967] <= 32'd8043;
		word[15'd8968] <= 32'd8044;
		word[15'd8969] <= 32'd8045;
		word[15'd8970] <= 32'd8046;
		word[15'd8971] <= 32'd8047;
		word[15'd8972] <= 32'd8048;
		word[15'd8973] <= 32'd8049;
		word[15'd8974] <= 32'd8050;
		word[15'd8975] <= 32'd8051;
		word[15'd8976] <= 32'd8052;
		word[15'd8977] <= 32'd8053;
		word[15'd8978] <= 32'd8054;
		word[15'd8979] <= 32'd8055;
		word[15'd8980] <= 32'd8056;
		word[15'd8981] <= 32'd8057;
		word[15'd8982] <= 32'd8058;
		word[15'd8983] <= 32'd8059;
		word[15'd8984] <= 32'd8060;
		word[15'd8985] <= 32'd8061;
		word[15'd8986] <= 32'd8062;
		word[15'd8987] <= 32'd8063;
		word[15'd8988] <= 32'd8064;
		word[15'd8989] <= 32'd8065;
		word[15'd8990] <= 32'd8066;
		word[15'd8991] <= 32'd8067;
		word[15'd8992] <= 32'd8068;
		word[15'd8993] <= 32'd8069;
		word[15'd8994] <= 32'd8070;
		word[15'd8995] <= 32'd8071;
		word[15'd8996] <= 32'd8072;
		word[15'd8997] <= 32'd8073;
		word[15'd8998] <= 32'd8074;
		word[15'd8999] <= 32'd8075;
		word[15'd9000] <= 32'd8076;
		word[15'd9001] <= 32'd8077;
		word[15'd9002] <= 32'd8078;
		word[15'd9003] <= 32'd8079;
		word[15'd9004] <= 32'd8080;
		word[15'd9005] <= 32'd8081;
		word[15'd9006] <= 32'd8082;
		word[15'd9007] <= 32'd8083;
		word[15'd9008] <= 32'd8084;
		word[15'd9009] <= 32'd8085;
		word[15'd9010] <= 32'd8086;
		word[15'd9011] <= 32'd8087;
		word[15'd9012] <= 32'd8088;
		word[15'd9013] <= 32'd8089;
		word[15'd9014] <= 32'd8090;
		word[15'd9015] <= 32'd8091;
		word[15'd9016] <= 32'd8092;
		word[15'd9017] <= 32'd8093;
		word[15'd9018] <= 32'd8094;
		word[15'd9019] <= 32'd8095;
		word[15'd9020] <= 32'd8096;
		word[15'd9021] <= 32'd8097;
		word[15'd9022] <= 32'd8098;
		word[15'd9023] <= 32'd8099;
		word[15'd9024] <= 32'd8100;
		word[15'd9025] <= 32'd8101;
		word[15'd9026] <= 32'd8102;
		word[15'd9027] <= 32'd8103;
		word[15'd9028] <= 32'd8104;
		word[15'd9029] <= 32'd8105;
		word[15'd9030] <= 32'd8106;
		word[15'd9031] <= 32'd8107;
		word[15'd9032] <= 32'd8108;
		word[15'd9033] <= 32'd8109;
		word[15'd9034] <= 32'd8110;
		word[15'd9035] <= 32'd8111;
		word[15'd9036] <= 32'd8112;
		word[15'd9037] <= 32'd8113;
		word[15'd9038] <= 32'd8114;
		word[15'd9039] <= 32'd8115;
		word[15'd9040] <= 32'd8116;
		word[15'd9041] <= 32'd8117;
		word[15'd9042] <= 32'd8118;
		word[15'd9043] <= 32'd8119;
		word[15'd9044] <= 32'd8120;
		word[15'd9045] <= 32'd8121;
		word[15'd9046] <= 32'd8122;
		word[15'd9047] <= 32'd8123;
		word[15'd9048] <= 32'd8124;
		word[15'd9049] <= 32'd8125;
		word[15'd9050] <= 32'd8126;
		word[15'd9051] <= 32'd8127;
		word[15'd9052] <= 32'd8128;
		word[15'd9053] <= 32'd8129;
		word[15'd9054] <= 32'd8130;
		word[15'd9055] <= 32'd8131;
		word[15'd9056] <= 32'd8132;
		word[15'd9057] <= 32'd8133;
		word[15'd9058] <= 32'd8134;
		word[15'd9059] <= 32'd8135;
		word[15'd9060] <= 32'd8136;
		word[15'd9061] <= 32'd8137;
		word[15'd9062] <= 32'd8138;
		word[15'd9063] <= 32'd8139;
		word[15'd9064] <= 32'd8140;
		word[15'd9065] <= 32'd8141;
		word[15'd9066] <= 32'd8142;
		word[15'd9067] <= 32'd8143;
		word[15'd9068] <= 32'd8144;
		word[15'd9069] <= 32'd8145;
		word[15'd9070] <= 32'd8146;
		word[15'd9071] <= 32'd8147;
		word[15'd9072] <= 32'd8148;
		word[15'd9073] <= 32'd8149;
		word[15'd9074] <= 32'd8150;
		word[15'd9075] <= 32'd8151;
		word[15'd9076] <= 32'd8152;
		word[15'd9077] <= 32'd8153;
		word[15'd9078] <= 32'd8154;
		word[15'd9079] <= 32'd8155;
		word[15'd9080] <= 32'd8156;
		word[15'd9081] <= 32'd8157;
		word[15'd9082] <= 32'd8158;
		word[15'd9083] <= 32'd8159;
		word[15'd9084] <= 32'd8160;
		word[15'd9085] <= 32'd8161;
		word[15'd9086] <= 32'd8162;
		word[15'd9087] <= 32'd8163;
		word[15'd9088] <= 32'd8164;
		word[15'd9089] <= 32'd8165;
		word[15'd9090] <= 32'd8166;
		word[15'd9091] <= 32'd8167;
		word[15'd9092] <= 32'd8168;
		word[15'd9093] <= 32'd8169;
		word[15'd9094] <= 32'd8170;
		word[15'd9095] <= 32'd8171;
		word[15'd9096] <= 32'd8172;
		word[15'd9097] <= 32'd8173;
		word[15'd9098] <= 32'd8174;
		word[15'd9099] <= 32'd8175;
		word[15'd9100] <= 32'd8176;
		word[15'd9101] <= 32'd8177;
		word[15'd9102] <= 32'd8178;
		word[15'd9103] <= 32'd8179;
		word[15'd9104] <= 32'd8180;
		word[15'd9105] <= 32'd8181;
		word[15'd9106] <= 32'd8182;
		word[15'd9107] <= 32'd8183;
		word[15'd9108] <= 32'd8184;
		word[15'd9109] <= 32'd8185;
		word[15'd9110] <= 32'd8186;
		word[15'd9111] <= 32'd8187;
		word[15'd9112] <= 32'd8188;
		word[15'd9113] <= 32'd8189;
		word[15'd9114] <= 32'd8190;
		word[15'd9115] <= 32'd8191;
		word[15'd9116] <= 32'd8192;
		word[15'd9117] <= 32'd8193;
		word[15'd9118] <= 32'd8194;
		word[15'd9119] <= 32'd8195;
		word[15'd9120] <= 32'd8196;
		word[15'd9121] <= 32'd8197;
		word[15'd9122] <= 32'd8198;
		word[15'd9123] <= 32'd8199;
		word[15'd9124] <= 32'd8200;
		word[15'd9125] <= 32'd8201;
		word[15'd9126] <= 32'd8202;
		word[15'd9127] <= 32'd8203;
		word[15'd9128] <= 32'd8204;
		word[15'd9129] <= 32'd8205;
		word[15'd9130] <= 32'd8206;
		word[15'd9131] <= 32'd8207;
		word[15'd9132] <= 32'd8208;
		word[15'd9133] <= 32'd8209;
		word[15'd9134] <= 32'd8210;
		word[15'd9135] <= 32'd8211;
		word[15'd9136] <= 32'd8212;
		word[15'd9137] <= 32'd8213;
		word[15'd9138] <= 32'd8214;
		word[15'd9139] <= 32'd8215;
		word[15'd9140] <= 32'd8216;
		word[15'd9141] <= 32'd8217;
		word[15'd9142] <= 32'd8218;
		word[15'd9143] <= 32'd8219;
		word[15'd9144] <= 32'd8220;
		word[15'd9145] <= 32'd8221;
		word[15'd9146] <= 32'd8222;
		word[15'd9147] <= 32'd8223;
		word[15'd9148] <= 32'd8224;
		word[15'd9149] <= 32'd8225;
		word[15'd9150] <= 32'd8226;
		word[15'd9151] <= 32'd8227;
		word[15'd9152] <= 32'd8228;
		word[15'd9153] <= 32'd8229;
		word[15'd9154] <= 32'd8230;
		word[15'd9155] <= 32'd8231;
		word[15'd9156] <= 32'd8232;
		word[15'd9157] <= 32'd8233;
		word[15'd9158] <= 32'd8234;
		word[15'd9159] <= 32'd8235;
		word[15'd9160] <= 32'd8236;
		word[15'd9161] <= 32'd8237;
		word[15'd9162] <= 32'd8238;
		word[15'd9163] <= 32'd8239;
		word[15'd9164] <= 32'd8240;
		word[15'd9165] <= 32'd8241;
		word[15'd9166] <= 32'd8242;
		word[15'd9167] <= 32'd8243;
		word[15'd9168] <= 32'd8244;
		word[15'd9169] <= 32'd8245;
		word[15'd9170] <= 32'd8246;
		word[15'd9171] <= 32'd8247;
		word[15'd9172] <= 32'd8248;
		word[15'd9173] <= 32'd8249;
		word[15'd9174] <= 32'd8250;
		word[15'd9175] <= 32'd8251;
		word[15'd9176] <= 32'd8252;
		word[15'd9177] <= 32'd8253;
		word[15'd9178] <= 32'd8254;
		word[15'd9179] <= 32'd8255;
		word[15'd9180] <= 32'd8256;
		word[15'd9181] <= 32'd8257;
		word[15'd9182] <= 32'd8258;
		word[15'd9183] <= 32'd8259;
		word[15'd9184] <= 32'd8260;
		word[15'd9185] <= 32'd8261;
		word[15'd9186] <= 32'd8262;
		word[15'd9187] <= 32'd8263;
		word[15'd9188] <= 32'd8264;
		word[15'd9189] <= 32'd8265;
		word[15'd9190] <= 32'd8266;
		word[15'd9191] <= 32'd8267;
		word[15'd9192] <= 32'd8268;
		word[15'd9193] <= 32'd8269;
		word[15'd9194] <= 32'd8270;
		word[15'd9195] <= 32'd8271;
		word[15'd9196] <= 32'd8272;
		word[15'd9197] <= 32'd8273;
		word[15'd9198] <= 32'd8274;
		word[15'd9199] <= 32'd8275;
		word[15'd9200] <= 32'd8276;
		word[15'd9201] <= 32'd8277;
		word[15'd9202] <= 32'd8278;
		word[15'd9203] <= 32'd8279;
		word[15'd9204] <= 32'd8280;
		word[15'd9205] <= 32'd8281;
		word[15'd9206] <= 32'd8282;
		word[15'd9207] <= 32'd8283;
		word[15'd9208] <= 32'd8284;
		word[15'd9209] <= 32'd8285;
		word[15'd9210] <= 32'd8286;
		word[15'd9211] <= 32'd8287;
		word[15'd9212] <= 32'd8288;
		word[15'd9213] <= 32'd8289;
		word[15'd9214] <= 32'd8290;
		word[15'd9215] <= 32'd8291;
		

	end



endmodule 